
module circuit ( CLK, RESET, DONE, MESSAGE1, MESSAGE2, MESSAGE3, RESULT1, 
        RESULT2, RESULT3 );
  input [199:0] MESSAGE1;
  input [199:0] MESSAGE2;
  input [199:0] MESSAGE3;
  output [199:0] RESULT1;
  output [199:0] RESULT2;
  output [199:0] RESULT3;
  input CLK, RESET;
  output DONE;
  wire   RoundFunction_T1_n600, RoundFunction_T1_n599, RoundFunction_T1_n598,
         RoundFunction_T1_n597, RoundFunction_T1_n596, RoundFunction_T1_n595,
         RoundFunction_T1_n594, RoundFunction_T1_n593, RoundFunction_T1_n592,
         RoundFunction_T1_n591, RoundFunction_T1_n590, RoundFunction_T1_n589,
         RoundFunction_T1_n588, RoundFunction_T1_n587, RoundFunction_T1_n586,
         RoundFunction_T1_n585, RoundFunction_T1_n584, RoundFunction_T1_n583,
         RoundFunction_T1_n582, RoundFunction_T1_n581, RoundFunction_T1_n580,
         RoundFunction_T1_n579, RoundFunction_T1_n578, RoundFunction_T1_n577,
         RoundFunction_T1_n576, RoundFunction_T1_n575, RoundFunction_T1_n574,
         RoundFunction_T1_n573, RoundFunction_T1_n572, RoundFunction_T1_n571,
         RoundFunction_T1_n570, RoundFunction_T1_n569, RoundFunction_T1_n568,
         RoundFunction_T1_n567, RoundFunction_T1_n566, RoundFunction_T1_n565,
         RoundFunction_T1_n564, RoundFunction_T1_n563, RoundFunction_T1_n562,
         RoundFunction_T1_n561, RoundFunction_T1_n560, RoundFunction_T1_n559,
         RoundFunction_T1_n558, RoundFunction_T1_n557, RoundFunction_T1_n556,
         RoundFunction_T1_n555, RoundFunction_T1_n554, RoundFunction_T1_n553,
         RoundFunction_T1_n552, RoundFunction_T1_n551, RoundFunction_T1_n550,
         RoundFunction_T1_n549, RoundFunction_T1_n548, RoundFunction_T1_n547,
         RoundFunction_T1_n546, RoundFunction_T1_n545, RoundFunction_T1_n544,
         RoundFunction_T1_n543, RoundFunction_T1_n542, RoundFunction_T1_n541,
         RoundFunction_T1_n540, RoundFunction_T1_n539, RoundFunction_T1_n538,
         RoundFunction_T1_n537, RoundFunction_T1_n536, RoundFunction_T1_n535,
         RoundFunction_T1_n534, RoundFunction_T1_n533, RoundFunction_T1_n532,
         RoundFunction_T1_n531, RoundFunction_T1_n530, RoundFunction_T1_n529,
         RoundFunction_T1_n528, RoundFunction_T1_n527, RoundFunction_T1_n526,
         RoundFunction_T1_n525, RoundFunction_T1_n524, RoundFunction_T1_n523,
         RoundFunction_T1_n522, RoundFunction_T1_n521, RoundFunction_T1_n520,
         RoundFunction_T1_n519, RoundFunction_T1_n518, RoundFunction_T1_n517,
         RoundFunction_T1_n516, RoundFunction_T1_n515, RoundFunction_T1_n514,
         RoundFunction_T1_n513, RoundFunction_T1_n512, RoundFunction_T1_n511,
         RoundFunction_T1_n510, RoundFunction_T1_n509, RoundFunction_T1_n508,
         RoundFunction_T1_n507, RoundFunction_T1_n506, RoundFunction_T1_n505,
         RoundFunction_T1_n504, RoundFunction_T1_n503, RoundFunction_T1_n502,
         RoundFunction_T1_n501, RoundFunction_T1_n500, RoundFunction_T1_n499,
         RoundFunction_T1_n498, RoundFunction_T1_n497, RoundFunction_T1_n496,
         RoundFunction_T1_n495, RoundFunction_T1_n494, RoundFunction_T1_n493,
         RoundFunction_T1_n492, RoundFunction_T1_n491, RoundFunction_T1_n490,
         RoundFunction_T1_n489, RoundFunction_T1_n488, RoundFunction_T1_n487,
         RoundFunction_T1_n486, RoundFunction_T1_n485, RoundFunction_T1_n484,
         RoundFunction_T1_n483, RoundFunction_T1_n482, RoundFunction_T1_n481,
         RoundFunction_T1_n480, RoundFunction_T1_n479, RoundFunction_T1_n478,
         RoundFunction_T1_n477, RoundFunction_T1_n476, RoundFunction_T1_n475,
         RoundFunction_T1_n474, RoundFunction_T1_n473, RoundFunction_T1_n472,
         RoundFunction_T1_n471, RoundFunction_T1_n470, RoundFunction_T1_n469,
         RoundFunction_T1_n468, RoundFunction_T1_n467, RoundFunction_T1_n466,
         RoundFunction_T1_n465, RoundFunction_T1_n464, RoundFunction_T1_n463,
         RoundFunction_T1_n462, RoundFunction_T1_n461, RoundFunction_T1_n460,
         RoundFunction_T1_n459, RoundFunction_T1_n458, RoundFunction_T1_n457,
         RoundFunction_T1_n456, RoundFunction_T1_n455, RoundFunction_T1_n454,
         RoundFunction_T1_n453, RoundFunction_T1_n452, RoundFunction_T1_n451,
         RoundFunction_T1_n450, RoundFunction_T1_n449, RoundFunction_T1_n448,
         RoundFunction_T1_n447, RoundFunction_T1_n446, RoundFunction_T1_n445,
         RoundFunction_T1_n444, RoundFunction_T1_n443, RoundFunction_T1_n442,
         RoundFunction_T1_n441, RoundFunction_T1_n440, RoundFunction_T1_n439,
         RoundFunction_T1_n438, RoundFunction_T1_n437, RoundFunction_T1_n436,
         RoundFunction_T1_n435, RoundFunction_T1_n434, RoundFunction_T1_n433,
         RoundFunction_T1_n432, RoundFunction_T1_n431, RoundFunction_T1_n430,
         RoundFunction_T1_n429, RoundFunction_T1_n428, RoundFunction_T1_n427,
         RoundFunction_T1_n426, RoundFunction_T1_n425, RoundFunction_T1_n424,
         RoundFunction_T1_n423, RoundFunction_T1_n422, RoundFunction_T1_n421,
         RoundFunction_T1_n420, RoundFunction_T1_n419, RoundFunction_T1_n418,
         RoundFunction_T1_n417, RoundFunction_T1_n416, RoundFunction_T1_n415,
         RoundFunction_T1_n414, RoundFunction_T1_n413, RoundFunction_T1_n412,
         RoundFunction_T1_n411, RoundFunction_T1_n410, RoundFunction_T1_n409,
         RoundFunction_T1_n408, RoundFunction_T1_n407, RoundFunction_T1_n406,
         RoundFunction_T1_n405, RoundFunction_T1_n404, RoundFunction_T1_n403,
         RoundFunction_T1_n402, RoundFunction_T1_n401, RoundFunction_T2_n600,
         RoundFunction_T2_n599, RoundFunction_T2_n598, RoundFunction_T2_n597,
         RoundFunction_T2_n596, RoundFunction_T2_n595, RoundFunction_T2_n594,
         RoundFunction_T2_n593, RoundFunction_T2_n592, RoundFunction_T2_n591,
         RoundFunction_T2_n590, RoundFunction_T2_n589, RoundFunction_T2_n588,
         RoundFunction_T2_n587, RoundFunction_T2_n586, RoundFunction_T2_n585,
         RoundFunction_T2_n584, RoundFunction_T2_n583, RoundFunction_T2_n582,
         RoundFunction_T2_n581, RoundFunction_T2_n580, RoundFunction_T2_n579,
         RoundFunction_T2_n578, RoundFunction_T2_n577, RoundFunction_T2_n576,
         RoundFunction_T2_n575, RoundFunction_T2_n574, RoundFunction_T2_n573,
         RoundFunction_T2_n572, RoundFunction_T2_n571, RoundFunction_T2_n570,
         RoundFunction_T2_n569, RoundFunction_T2_n568, RoundFunction_T2_n567,
         RoundFunction_T2_n566, RoundFunction_T2_n565, RoundFunction_T2_n564,
         RoundFunction_T2_n563, RoundFunction_T2_n562, RoundFunction_T2_n561,
         RoundFunction_T2_n560, RoundFunction_T2_n559, RoundFunction_T2_n558,
         RoundFunction_T2_n557, RoundFunction_T2_n556, RoundFunction_T2_n555,
         RoundFunction_T2_n554, RoundFunction_T2_n553, RoundFunction_T2_n552,
         RoundFunction_T2_n551, RoundFunction_T2_n550, RoundFunction_T2_n549,
         RoundFunction_T2_n548, RoundFunction_T2_n547, RoundFunction_T2_n546,
         RoundFunction_T2_n545, RoundFunction_T2_n544, RoundFunction_T2_n543,
         RoundFunction_T2_n542, RoundFunction_T2_n541, RoundFunction_T2_n540,
         RoundFunction_T2_n539, RoundFunction_T2_n538, RoundFunction_T2_n537,
         RoundFunction_T2_n536, RoundFunction_T2_n535, RoundFunction_T2_n534,
         RoundFunction_T2_n533, RoundFunction_T2_n532, RoundFunction_T2_n531,
         RoundFunction_T2_n530, RoundFunction_T2_n529, RoundFunction_T2_n528,
         RoundFunction_T2_n527, RoundFunction_T2_n526, RoundFunction_T2_n525,
         RoundFunction_T2_n524, RoundFunction_T2_n523, RoundFunction_T2_n522,
         RoundFunction_T2_n521, RoundFunction_T2_n520, RoundFunction_T2_n519,
         RoundFunction_T2_n518, RoundFunction_T2_n517, RoundFunction_T2_n516,
         RoundFunction_T2_n515, RoundFunction_T2_n514, RoundFunction_T2_n513,
         RoundFunction_T2_n512, RoundFunction_T2_n511, RoundFunction_T2_n510,
         RoundFunction_T2_n509, RoundFunction_T2_n508, RoundFunction_T2_n507,
         RoundFunction_T2_n506, RoundFunction_T2_n505, RoundFunction_T2_n504,
         RoundFunction_T2_n503, RoundFunction_T2_n502, RoundFunction_T2_n501,
         RoundFunction_T2_n500, RoundFunction_T2_n499, RoundFunction_T2_n498,
         RoundFunction_T2_n497, RoundFunction_T2_n496, RoundFunction_T2_n495,
         RoundFunction_T2_n494, RoundFunction_T2_n493, RoundFunction_T2_n492,
         RoundFunction_T2_n491, RoundFunction_T2_n490, RoundFunction_T2_n489,
         RoundFunction_T2_n488, RoundFunction_T2_n487, RoundFunction_T2_n486,
         RoundFunction_T2_n485, RoundFunction_T2_n484, RoundFunction_T2_n483,
         RoundFunction_T2_n482, RoundFunction_T2_n481, RoundFunction_T2_n480,
         RoundFunction_T2_n479, RoundFunction_T2_n478, RoundFunction_T2_n477,
         RoundFunction_T2_n476, RoundFunction_T2_n475, RoundFunction_T2_n474,
         RoundFunction_T2_n473, RoundFunction_T2_n472, RoundFunction_T2_n471,
         RoundFunction_T2_n470, RoundFunction_T2_n469, RoundFunction_T2_n468,
         RoundFunction_T2_n467, RoundFunction_T2_n466, RoundFunction_T2_n465,
         RoundFunction_T2_n464, RoundFunction_T2_n463, RoundFunction_T2_n462,
         RoundFunction_T2_n461, RoundFunction_T2_n460, RoundFunction_T2_n459,
         RoundFunction_T2_n458, RoundFunction_T2_n457, RoundFunction_T2_n456,
         RoundFunction_T2_n455, RoundFunction_T2_n454, RoundFunction_T2_n453,
         RoundFunction_T2_n452, RoundFunction_T2_n451, RoundFunction_T2_n450,
         RoundFunction_T2_n449, RoundFunction_T2_n448, RoundFunction_T2_n447,
         RoundFunction_T2_n446, RoundFunction_T2_n445, RoundFunction_T2_n444,
         RoundFunction_T2_n443, RoundFunction_T2_n442, RoundFunction_T2_n441,
         RoundFunction_T2_n440, RoundFunction_T2_n439, RoundFunction_T2_n438,
         RoundFunction_T2_n437, RoundFunction_T2_n436, RoundFunction_T2_n435,
         RoundFunction_T2_n434, RoundFunction_T2_n433, RoundFunction_T2_n432,
         RoundFunction_T2_n431, RoundFunction_T2_n430, RoundFunction_T2_n429,
         RoundFunction_T2_n428, RoundFunction_T2_n427, RoundFunction_T2_n426,
         RoundFunction_T2_n425, RoundFunction_T2_n424, RoundFunction_T2_n423,
         RoundFunction_T2_n422, RoundFunction_T2_n421, RoundFunction_T2_n420,
         RoundFunction_T2_n419, RoundFunction_T2_n418, RoundFunction_T2_n417,
         RoundFunction_T2_n416, RoundFunction_T2_n415, RoundFunction_T2_n414,
         RoundFunction_T2_n413, RoundFunction_T2_n412, RoundFunction_T2_n411,
         RoundFunction_T2_n410, RoundFunction_T2_n409, RoundFunction_T2_n408,
         RoundFunction_T2_n407, RoundFunction_T2_n406, RoundFunction_T2_n405,
         RoundFunction_T2_n404, RoundFunction_T2_n403, RoundFunction_T2_n402,
         RoundFunction_T2_n401, RoundFunction_T3_n600, RoundFunction_T3_n599,
         RoundFunction_T3_n598, RoundFunction_T3_n597, RoundFunction_T3_n596,
         RoundFunction_T3_n595, RoundFunction_T3_n594, RoundFunction_T3_n593,
         RoundFunction_T3_n592, RoundFunction_T3_n591, RoundFunction_T3_n590,
         RoundFunction_T3_n589, RoundFunction_T3_n588, RoundFunction_T3_n587,
         RoundFunction_T3_n586, RoundFunction_T3_n585, RoundFunction_T3_n584,
         RoundFunction_T3_n583, RoundFunction_T3_n582, RoundFunction_T3_n581,
         RoundFunction_T3_n580, RoundFunction_T3_n579, RoundFunction_T3_n578,
         RoundFunction_T3_n577, RoundFunction_T3_n576, RoundFunction_T3_n575,
         RoundFunction_T3_n574, RoundFunction_T3_n573, RoundFunction_T3_n572,
         RoundFunction_T3_n571, RoundFunction_T3_n570, RoundFunction_T3_n569,
         RoundFunction_T3_n568, RoundFunction_T3_n567, RoundFunction_T3_n566,
         RoundFunction_T3_n565, RoundFunction_T3_n564, RoundFunction_T3_n563,
         RoundFunction_T3_n562, RoundFunction_T3_n561, RoundFunction_T3_n560,
         RoundFunction_T3_n559, RoundFunction_T3_n558, RoundFunction_T3_n557,
         RoundFunction_T3_n556, RoundFunction_T3_n555, RoundFunction_T3_n554,
         RoundFunction_T3_n553, RoundFunction_T3_n552, RoundFunction_T3_n551,
         RoundFunction_T3_n550, RoundFunction_T3_n549, RoundFunction_T3_n548,
         RoundFunction_T3_n547, RoundFunction_T3_n546, RoundFunction_T3_n545,
         RoundFunction_T3_n544, RoundFunction_T3_n543, RoundFunction_T3_n542,
         RoundFunction_T3_n541, RoundFunction_T3_n540, RoundFunction_T3_n539,
         RoundFunction_T3_n538, RoundFunction_T3_n537, RoundFunction_T3_n536,
         RoundFunction_T3_n535, RoundFunction_T3_n534, RoundFunction_T3_n533,
         RoundFunction_T3_n532, RoundFunction_T3_n531, RoundFunction_T3_n530,
         RoundFunction_T3_n529, RoundFunction_T3_n528, RoundFunction_T3_n527,
         RoundFunction_T3_n526, RoundFunction_T3_n525, RoundFunction_T3_n524,
         RoundFunction_T3_n523, RoundFunction_T3_n522, RoundFunction_T3_n521,
         RoundFunction_T3_n520, RoundFunction_T3_n519, RoundFunction_T3_n518,
         RoundFunction_T3_n517, RoundFunction_T3_n516, RoundFunction_T3_n515,
         RoundFunction_T3_n514, RoundFunction_T3_n513, RoundFunction_T3_n512,
         RoundFunction_T3_n511, RoundFunction_T3_n510, RoundFunction_T3_n509,
         RoundFunction_T3_n508, RoundFunction_T3_n507, RoundFunction_T3_n506,
         RoundFunction_T3_n505, RoundFunction_T3_n504, RoundFunction_T3_n503,
         RoundFunction_T3_n502, RoundFunction_T3_n501, RoundFunction_T3_n500,
         RoundFunction_T3_n499, RoundFunction_T3_n498, RoundFunction_T3_n497,
         RoundFunction_T3_n496, RoundFunction_T3_n495, RoundFunction_T3_n494,
         RoundFunction_T3_n493, RoundFunction_T3_n492, RoundFunction_T3_n491,
         RoundFunction_T3_n490, RoundFunction_T3_n489, RoundFunction_T3_n488,
         RoundFunction_T3_n487, RoundFunction_T3_n486, RoundFunction_T3_n485,
         RoundFunction_T3_n484, RoundFunction_T3_n483, RoundFunction_T3_n482,
         RoundFunction_T3_n481, RoundFunction_T3_n480, RoundFunction_T3_n479,
         RoundFunction_T3_n478, RoundFunction_T3_n477, RoundFunction_T3_n476,
         RoundFunction_T3_n475, RoundFunction_T3_n474, RoundFunction_T3_n473,
         RoundFunction_T3_n472, RoundFunction_T3_n471, RoundFunction_T3_n470,
         RoundFunction_T3_n469, RoundFunction_T3_n468, RoundFunction_T3_n467,
         RoundFunction_T3_n466, RoundFunction_T3_n465, RoundFunction_T3_n464,
         RoundFunction_T3_n463, RoundFunction_T3_n462, RoundFunction_T3_n461,
         RoundFunction_T3_n460, RoundFunction_T3_n459, RoundFunction_T3_n458,
         RoundFunction_T3_n457, RoundFunction_T3_n456, RoundFunction_T3_n455,
         RoundFunction_T3_n454, RoundFunction_T3_n453, RoundFunction_T3_n452,
         RoundFunction_T3_n451, RoundFunction_T3_n450, RoundFunction_T3_n449,
         RoundFunction_T3_n448, RoundFunction_T3_n447, RoundFunction_T3_n446,
         RoundFunction_T3_n445, RoundFunction_T3_n444, RoundFunction_T3_n443,
         RoundFunction_T3_n442, RoundFunction_T3_n441, RoundFunction_T3_n440,
         RoundFunction_T3_n439, RoundFunction_T3_n438, RoundFunction_T3_n437,
         RoundFunction_T3_n436, RoundFunction_T3_n435, RoundFunction_T3_n434,
         RoundFunction_T3_n433, RoundFunction_T3_n432, RoundFunction_T3_n431,
         RoundFunction_T3_n430, RoundFunction_T3_n429, RoundFunction_T3_n428,
         RoundFunction_T3_n427, RoundFunction_T3_n426, RoundFunction_T3_n425,
         RoundFunction_T3_n424, RoundFunction_T3_n423, RoundFunction_T3_n422,
         RoundFunction_T3_n421, RoundFunction_T3_n420, RoundFunction_T3_n419,
         RoundFunction_T3_n418, RoundFunction_T3_n417, RoundFunction_T3_n416,
         RoundFunction_T3_n415, RoundFunction_T3_n414, RoundFunction_T3_n413,
         RoundFunction_T3_n412, RoundFunction_T3_n411, RoundFunction_T3_n410,
         RoundFunction_T3_n409, RoundFunction_T3_n408, RoundFunction_T3_n407,
         RoundFunction_T3_n406, RoundFunction_T3_n405, RoundFunction_T3_n404,
         RoundFunction_T3_n403, RoundFunction_T3_n402, RoundFunction_T3_n401,
         RoundFunction_C_Inst_Chi_NoFresh_0_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_0_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_0_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_0_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_0_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_0_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_0_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_0_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_0_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_0_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_0_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_0_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_0_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_0_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_0_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_1_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_1_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_1_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_1_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_1_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_1_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_1_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_1_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_1_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_1_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_1_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_1_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_1_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_1_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_2_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_2_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_2_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_2_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_2_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_2_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_2_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_2_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_2_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_2_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_2_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_2_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_2_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_2_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_3_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_3_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_3_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_3_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_3_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_3_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_3_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_3_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_3_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_3_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_3_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_3_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_3_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_3_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_4_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_4_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_4_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_4_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_4_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_4_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_4_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_4_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_4_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_4_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_4_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_4_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_4_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_4_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_5_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_5_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_5_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_5_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_5_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_5_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_5_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_5_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_5_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_5_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_5_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_5_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_5_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_5_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_6_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_6_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_6_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_6_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_6_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_6_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_6_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_6_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_6_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_6_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_6_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_6_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_6_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_6_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_7_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_7_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_7_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_7_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_7_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_7_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_7_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_7_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_7_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_7_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_7_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_7_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_7_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_7_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_8_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_8_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_8_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_8_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_8_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_8_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_8_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_8_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_8_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_8_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_8_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_8_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_8_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_8_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_9_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_9_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_9_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_9_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_9_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_9_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_9_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_9_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_9_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_9_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_9_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_9_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_9_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_9_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_10_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_10_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_10_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_10_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_10_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_10_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_10_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_10_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_10_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_10_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_10_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_10_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_10_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_10_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_11_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_11_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_11_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_11_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_11_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_11_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_11_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_11_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_11_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_11_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_11_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_11_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_11_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_11_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_12_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_12_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_12_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_12_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_12_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_12_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_12_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_12_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_12_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_12_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_12_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_12_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_12_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_12_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_13_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_13_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_13_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_13_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_13_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_13_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_13_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_13_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_13_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_13_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_13_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_13_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_13_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_13_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_14_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_14_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_14_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_14_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_14_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_14_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_14_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_14_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_14_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_14_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_14_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_14_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_14_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_14_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_15_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_15_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_15_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_15_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_15_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_15_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_15_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_15_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_15_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_15_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_15_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_15_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_15_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_15_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_16_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_16_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_16_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_16_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_16_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_16_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_16_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_16_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_16_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_16_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_16_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_16_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_16_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_16_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_17_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_17_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_17_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_17_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_17_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_17_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_17_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_17_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_17_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_17_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_17_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_17_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_17_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_17_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_18_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_18_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_18_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_18_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_18_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_18_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_18_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_18_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_18_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_18_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_18_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_18_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_18_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_18_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_19_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_19_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_19_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_19_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_19_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_19_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_19_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_19_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_19_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_19_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_19_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_19_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_19_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_19_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_20_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_20_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_20_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_20_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_20_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_20_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_20_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_20_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_20_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_20_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_20_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_20_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_20_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_20_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_21_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_21_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_21_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_21_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_21_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_21_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_21_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_21_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_21_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_21_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_21_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_21_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_21_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_21_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_22_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_22_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_22_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_22_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_22_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_22_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_22_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_22_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_22_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_22_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_22_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_22_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_22_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_22_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_23_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_23_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_23_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_23_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_23_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_23_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_23_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_23_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_23_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_23_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_23_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_23_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_23_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_23_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_24_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_24_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_24_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_24_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_24_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_24_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_24_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_24_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_24_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_24_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_24_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_24_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_24_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_24_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_25_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_25_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_25_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_25_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_25_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_25_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_25_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_25_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_25_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_25_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_25_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_25_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_25_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_25_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_26_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_26_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_26_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_26_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_26_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_26_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_26_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_26_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_26_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_26_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_26_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_26_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_26_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_26_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_27_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_27_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_27_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_27_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_27_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_27_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_27_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_27_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_27_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_27_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_27_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_27_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_27_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_27_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_28_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_28_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_28_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_28_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_28_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_28_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_28_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_28_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_28_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_28_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_28_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_28_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_28_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_28_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_29_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_29_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_29_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_29_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_29_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_29_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_29_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_29_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_29_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_29_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_29_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_29_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_29_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_29_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_30_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_30_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_30_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_30_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_30_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_30_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_30_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_30_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_30_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_30_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_30_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_30_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_30_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_30_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_31_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_31_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_31_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_31_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_31_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_31_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_31_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_31_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_31_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_31_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_31_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_31_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_31_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_31_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_32_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_32_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_32_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_32_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_32_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_32_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_32_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_32_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_32_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_32_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_32_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_32_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_32_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_32_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_33_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_33_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_33_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_33_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_33_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_33_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_33_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_33_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_33_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_33_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_33_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_33_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_33_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_33_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_34_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_34_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_34_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_34_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_34_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_34_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_34_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_34_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_34_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_34_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_34_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_34_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_34_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_34_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_35_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_35_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_35_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_35_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_35_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_35_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_35_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_35_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_35_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_35_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_35_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_35_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_35_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_35_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_36_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_36_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_36_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_36_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_36_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_36_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_36_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_36_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_36_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_36_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_36_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_36_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_36_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_36_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_37_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_37_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_37_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_37_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_37_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_37_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_37_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_37_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_37_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_37_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_37_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_37_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_37_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_37_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_38_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_38_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_38_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_38_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_38_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_38_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_38_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_38_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_38_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_38_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_38_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_38_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_38_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_38_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_e_1_,
         RoundFunction_C_Inst_Chi_NoFresh_39_e_2_,
         RoundFunction_C_Inst_Chi_NoFresh_39_e_3_,
         RoundFunction_C_Inst_Chi_NoFresh_39_d_1_,
         RoundFunction_C_Inst_Chi_NoFresh_39_d_2_,
         RoundFunction_C_Inst_Chi_NoFresh_39_d_3_,
         RoundFunction_C_Inst_Chi_NoFresh_39_c_1_,
         RoundFunction_C_Inst_Chi_NoFresh_39_c_2_,
         RoundFunction_C_Inst_Chi_NoFresh_39_c_3_,
         RoundFunction_C_Inst_Chi_NoFresh_39_b_1_,
         RoundFunction_C_Inst_Chi_NoFresh_39_b_2_,
         RoundFunction_C_Inst_Chi_NoFresh_39_b_3_,
         RoundFunction_C_Inst_Chi_NoFresh_39_a_1_,
         RoundFunction_C_Inst_Chi_NoFresh_39_a_2_,
         RoundFunction_C_Inst_Chi_NoFresh_39_a_3_,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_1__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_3__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_5__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_6__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_8__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_8__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_9__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_10__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_11__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_12__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_14__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_14__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_15__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_17__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_20__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_21__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_23__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_24__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_24__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_25__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_29__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_29__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_30__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_32__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_32__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_33__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_34__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_35__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_38__CF_Inst_n7,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_39__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_41__CF_Inst_n6,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_41__CF_Inst_n5,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_42__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_Inst_44__CF_Inst_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression3_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression1_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression2_n3,
         RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression3_n3,
         FSM_n92, FSM_n91, FSM_n90, FSM_n89, FSM_n88, FSM_n86, FSM_n85,
         FSM_n84, FSM_n83, FSM_n82, FSM_n81, FSM_n80, FSM_n69, FSM_n68,
         FSM_n67, FSM_n66, FSM_n65, FSM_n64, FSM_n63, FSM_n62, FSM_n61,
         FSM_n60, FSM_n59, FSM_n58, FSM_n57, FSM_n56, FSM_n55, FSM_n54,
         FSM_n53, FSM_n52, FSM_n51, FSM_n50, FSM_n49, FSM_n48, FSM_n47,
         FSM_n46, FSM_n45, FSM_n44, FSM_n43, FSM_n42, FSM_n41, FSM_n40,
         FSM_n39, FSM_n38, FSM_n37, FSM_n36, FSM_n35, FSM_n34, FSM_n33,
         FSM_n32, FSM_n31, FSM_n30, FSM_n29, FSM_n28, FSM_n27, FSM_n26,
         FSM_n25, FSM_n24, FSM_n23, FSM_n22, FSM_n21, FSM_n20, FSM_n87, FSM_n1,
         FSM_n79, FSM_n78, FSM_n77, FSM_n76, FSM_n75, FSM_n74, FSM_n73,
         FSM_n72, FSM_n71, FSM_n70, FSM_n18, FSM_n17, FSM_n15, FSM_n14,
         FSM_n13, FSM_n12, FSM_n11, FSM_n10, FSM_n8, FSM_n7,
         FSM_CONST_internal_3, FSM_CONST_internal_7;
  wire   [7:0] CONST;
  wire   [199:0] RoundFunction_TMP3_3;
  wire   [199:0] RoundFunction_TMP3_2;
  wire   [7:0] RoundFunction_TMP4_1;
  wire   [199:0] RoundFunction_TMP3_1;
  wire   [199:0] RoundFunction_STATE3;
  wire   [199:0] RoundFunction_STATE2;
  wire   [199:0] RoundFunction_STATE1;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg;
  wire   [44:0] RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out;
  wire   [1:0] FSM_CONST_internal;

  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_0_ ( .D(RESULT1[192]), 
        .SI(MESSAGE1[192]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[0]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_1_ ( .D(RESULT1[193]), 
        .SI(MESSAGE1[193]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[1]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_2_ ( .D(RESULT1[194]), 
        .SI(MESSAGE1[194]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[2]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_3_ ( .D(RESULT1[195]), 
        .SI(MESSAGE1[195]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[3]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_4_ ( .D(RESULT1[196]), 
        .SI(MESSAGE1[196]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[4]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_5_ ( .D(RESULT1[197]), 
        .SI(MESSAGE1[197]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[5]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_6_ ( .D(RESULT1[198]), 
        .SI(MESSAGE1[198]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[6]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_7_ ( .D(RESULT1[199]), 
        .SI(MESSAGE1[199]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[7]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_8_ ( .D(RESULT1[184]), 
        .SI(MESSAGE1[184]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[8]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_9_ ( .D(RESULT1[185]), 
        .SI(MESSAGE1[185]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[9]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_10_ ( .D(RESULT1[186]), 
        .SI(MESSAGE1[186]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[10]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_11_ ( .D(RESULT1[187]), 
        .SI(MESSAGE1[187]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[11]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_12_ ( .D(RESULT1[188]), 
        .SI(MESSAGE1[188]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[12]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_13_ ( .D(RESULT1[189]), 
        .SI(MESSAGE1[189]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[13]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_14_ ( .D(RESULT1[190]), 
        .SI(MESSAGE1[190]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[14]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_15_ ( .D(RESULT1[191]), 
        .SI(MESSAGE1[191]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[15]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_16_ ( .D(RESULT1[176]), 
        .SI(MESSAGE1[176]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[16]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_17_ ( .D(RESULT1[177]), 
        .SI(MESSAGE1[177]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[17]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_18_ ( .D(RESULT1[178]), 
        .SI(MESSAGE1[178]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[18]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_19_ ( .D(RESULT1[179]), 
        .SI(MESSAGE1[179]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[19]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_20_ ( .D(RESULT1[180]), 
        .SI(MESSAGE1[180]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[20]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_21_ ( .D(RESULT1[181]), 
        .SI(MESSAGE1[181]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[21]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_22_ ( .D(RESULT1[182]), 
        .SI(MESSAGE1[182]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[22]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_23_ ( .D(RESULT1[183]), 
        .SI(MESSAGE1[183]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[23]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_24_ ( .D(RESULT1[168]), 
        .SI(MESSAGE1[168]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[24]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_25_ ( .D(RESULT1[169]), 
        .SI(MESSAGE1[169]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[25]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_26_ ( .D(RESULT1[170]), 
        .SI(MESSAGE1[170]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[26]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_27_ ( .D(RESULT1[171]), 
        .SI(MESSAGE1[171]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[27]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_28_ ( .D(RESULT1[172]), 
        .SI(MESSAGE1[172]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[28]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_29_ ( .D(RESULT1[173]), 
        .SI(MESSAGE1[173]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[29]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_30_ ( .D(RESULT1[174]), 
        .SI(MESSAGE1[174]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[30]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_31_ ( .D(RESULT1[175]), 
        .SI(MESSAGE1[175]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[31]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_32_ ( .D(RESULT1[160]), 
        .SI(MESSAGE1[160]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[32]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_33_ ( .D(RESULT1[161]), 
        .SI(MESSAGE1[161]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[33]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_34_ ( .D(RESULT1[162]), 
        .SI(MESSAGE1[162]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[34]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_35_ ( .D(RESULT1[163]), 
        .SI(MESSAGE1[163]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[35]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_36_ ( .D(RESULT1[164]), 
        .SI(MESSAGE1[164]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[36]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_37_ ( .D(RESULT1[165]), 
        .SI(MESSAGE1[165]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[37]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_38_ ( .D(RESULT1[166]), 
        .SI(MESSAGE1[166]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[38]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_39_ ( .D(RESULT1[167]), 
        .SI(MESSAGE1[167]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[39]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_40_ ( .D(RESULT1[152]), 
        .SI(MESSAGE1[152]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[40]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_41_ ( .D(RESULT1[153]), 
        .SI(MESSAGE1[153]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[41]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_42_ ( .D(RESULT1[154]), 
        .SI(MESSAGE1[154]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[42]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_43_ ( .D(RESULT1[155]), 
        .SI(MESSAGE1[155]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[43]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_44_ ( .D(RESULT1[156]), 
        .SI(MESSAGE1[156]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[44]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_45_ ( .D(RESULT1[157]), 
        .SI(MESSAGE1[157]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[45]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_46_ ( .D(RESULT1[158]), 
        .SI(MESSAGE1[158]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[46]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_47_ ( .D(RESULT1[159]), 
        .SI(MESSAGE1[159]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[47]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_48_ ( .D(RESULT1[144]), 
        .SI(MESSAGE1[144]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[48]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_49_ ( .D(RESULT1[145]), 
        .SI(MESSAGE1[145]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[49]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_50_ ( .D(RESULT1[146]), 
        .SI(MESSAGE1[146]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[50]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_51_ ( .D(RESULT1[147]), 
        .SI(MESSAGE1[147]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[51]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_52_ ( .D(RESULT1[148]), 
        .SI(MESSAGE1[148]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[52]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_53_ ( .D(RESULT1[149]), 
        .SI(MESSAGE1[149]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[53]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_54_ ( .D(RESULT1[150]), 
        .SI(MESSAGE1[150]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[54]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_55_ ( .D(RESULT1[151]), 
        .SI(MESSAGE1[151]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[55]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_56_ ( .D(RESULT1[136]), 
        .SI(MESSAGE1[136]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[56]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_57_ ( .D(RESULT1[137]), 
        .SI(MESSAGE1[137]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[57]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_58_ ( .D(RESULT1[138]), 
        .SI(MESSAGE1[138]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[58]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_59_ ( .D(RESULT1[139]), 
        .SI(MESSAGE1[139]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[59]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_60_ ( .D(RESULT1[140]), 
        .SI(MESSAGE1[140]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[60]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_61_ ( .D(RESULT1[141]), 
        .SI(MESSAGE1[141]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[61]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_62_ ( .D(RESULT1[142]), 
        .SI(MESSAGE1[142]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[62]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_63_ ( .D(RESULT1[143]), 
        .SI(MESSAGE1[143]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[63]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_64_ ( .D(RESULT1[128]), 
        .SI(MESSAGE1[128]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[64]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_65_ ( .D(RESULT1[129]), 
        .SI(MESSAGE1[129]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[65]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_66_ ( .D(RESULT1[130]), 
        .SI(MESSAGE1[130]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[66]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_67_ ( .D(RESULT1[131]), 
        .SI(MESSAGE1[131]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[67]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_68_ ( .D(RESULT1[132]), 
        .SI(MESSAGE1[132]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[68]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_69_ ( .D(RESULT1[133]), 
        .SI(MESSAGE1[133]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[69]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_70_ ( .D(RESULT1[134]), 
        .SI(MESSAGE1[134]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[70]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_71_ ( .D(RESULT1[135]), 
        .SI(MESSAGE1[135]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[71]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_72_ ( .D(RESULT1[120]), 
        .SI(MESSAGE1[120]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[72]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_73_ ( .D(RESULT1[121]), 
        .SI(MESSAGE1[121]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[73]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_74_ ( .D(RESULT1[122]), 
        .SI(MESSAGE1[122]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[74]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_75_ ( .D(RESULT1[123]), 
        .SI(MESSAGE1[123]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[75]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_76_ ( .D(RESULT1[124]), 
        .SI(MESSAGE1[124]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[76]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_77_ ( .D(RESULT1[125]), 
        .SI(MESSAGE1[125]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[77]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_78_ ( .D(RESULT1[126]), 
        .SI(MESSAGE1[126]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[78]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_79_ ( .D(RESULT1[127]), 
        .SI(MESSAGE1[127]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[79]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_80_ ( .D(RESULT1[112]), 
        .SI(MESSAGE1[112]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[80]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_81_ ( .D(RESULT1[113]), 
        .SI(MESSAGE1[113]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[81]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_82_ ( .D(RESULT1[114]), 
        .SI(MESSAGE1[114]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[82]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_83_ ( .D(RESULT1[115]), 
        .SI(MESSAGE1[115]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[83]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_84_ ( .D(RESULT1[116]), 
        .SI(MESSAGE1[116]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[84]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_85_ ( .D(RESULT1[117]), 
        .SI(MESSAGE1[117]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[85]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_86_ ( .D(RESULT1[118]), 
        .SI(MESSAGE1[118]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[86]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_87_ ( .D(RESULT1[119]), 
        .SI(MESSAGE1[119]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[87]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_88_ ( .D(RESULT1[104]), 
        .SI(MESSAGE1[104]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[88]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_89_ ( .D(RESULT1[105]), 
        .SI(MESSAGE1[105]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[89]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_90_ ( .D(RESULT1[106]), 
        .SI(MESSAGE1[106]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[90]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_91_ ( .D(RESULT1[107]), 
        .SI(MESSAGE1[107]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[91]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_92_ ( .D(RESULT1[108]), 
        .SI(MESSAGE1[108]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[92]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_93_ ( .D(RESULT1[109]), 
        .SI(MESSAGE1[109]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[93]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_94_ ( .D(RESULT1[110]), 
        .SI(MESSAGE1[110]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[94]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_95_ ( .D(RESULT1[111]), 
        .SI(MESSAGE1[111]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[95]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_96_ ( .D(RESULT1[96]), 
        .SI(MESSAGE1[96]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[96]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_97_ ( .D(RESULT1[97]), 
        .SI(MESSAGE1[97]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[97]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_98_ ( .D(RESULT1[98]), 
        .SI(MESSAGE1[98]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[98]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_99_ ( .D(RESULT1[99]), 
        .SI(MESSAGE1[99]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[99]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_100_ ( .D(RESULT1[100]), 
        .SI(MESSAGE1[100]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[100]), .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_101_ ( .D(RESULT1[101]), 
        .SI(MESSAGE1[101]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[101]), .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_102_ ( .D(RESULT1[102]), 
        .SI(MESSAGE1[102]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[102]), .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_103_ ( .D(RESULT1[103]), 
        .SI(MESSAGE1[103]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[103]), .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_104_ ( .D(RESULT1[88]), 
        .SI(MESSAGE1[88]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[104]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_105_ ( .D(RESULT1[89]), 
        .SI(MESSAGE1[89]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[105]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_106_ ( .D(RESULT1[90]), 
        .SI(MESSAGE1[90]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[106]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_107_ ( .D(RESULT1[91]), 
        .SI(MESSAGE1[91]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[107]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_108_ ( .D(RESULT1[92]), 
        .SI(MESSAGE1[92]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[108]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_109_ ( .D(RESULT1[93]), 
        .SI(MESSAGE1[93]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[109]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_110_ ( .D(RESULT1[94]), 
        .SI(MESSAGE1[94]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[110]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_111_ ( .D(RESULT1[95]), 
        .SI(MESSAGE1[95]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[111]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_112_ ( .D(RESULT1[80]), 
        .SI(MESSAGE1[80]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[112]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_113_ ( .D(RESULT1[81]), 
        .SI(MESSAGE1[81]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[113]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_114_ ( .D(RESULT1[82]), 
        .SI(MESSAGE1[82]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[114]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_115_ ( .D(RESULT1[83]), 
        .SI(MESSAGE1[83]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[115]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_116_ ( .D(RESULT1[84]), 
        .SI(MESSAGE1[84]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[116]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_117_ ( .D(RESULT1[85]), 
        .SI(MESSAGE1[85]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[117]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_118_ ( .D(RESULT1[86]), 
        .SI(MESSAGE1[86]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[118]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_119_ ( .D(RESULT1[87]), 
        .SI(MESSAGE1[87]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[119]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_120_ ( .D(RESULT1[72]), 
        .SI(MESSAGE1[72]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[120]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_121_ ( .D(RESULT1[73]), 
        .SI(MESSAGE1[73]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[121]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_122_ ( .D(RESULT1[74]), 
        .SI(MESSAGE1[74]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[122]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_123_ ( .D(RESULT1[75]), 
        .SI(MESSAGE1[75]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[123]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_124_ ( .D(RESULT1[76]), 
        .SI(MESSAGE1[76]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[124]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_125_ ( .D(RESULT1[77]), 
        .SI(MESSAGE1[77]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[125]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_126_ ( .D(RESULT1[78]), 
        .SI(MESSAGE1[78]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[126]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_127_ ( .D(RESULT1[79]), 
        .SI(MESSAGE1[79]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[127]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_128_ ( .D(RESULT1[64]), 
        .SI(MESSAGE1[64]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[128]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_129_ ( .D(RESULT1[65]), 
        .SI(MESSAGE1[65]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[129]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_130_ ( .D(RESULT1[66]), 
        .SI(MESSAGE1[66]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[130]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_131_ ( .D(RESULT1[67]), 
        .SI(MESSAGE1[67]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[131]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_132_ ( .D(RESULT1[68]), 
        .SI(MESSAGE1[68]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[132]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_133_ ( .D(RESULT1[69]), 
        .SI(MESSAGE1[69]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[133]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_134_ ( .D(RESULT1[70]), 
        .SI(MESSAGE1[70]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[134]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_135_ ( .D(RESULT1[71]), 
        .SI(MESSAGE1[71]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[135]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_136_ ( .D(RESULT1[56]), 
        .SI(MESSAGE1[56]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[136]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_137_ ( .D(RESULT1[57]), 
        .SI(MESSAGE1[57]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[137]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_138_ ( .D(RESULT1[58]), 
        .SI(MESSAGE1[58]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[138]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_139_ ( .D(RESULT1[59]), 
        .SI(MESSAGE1[59]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[139]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_140_ ( .D(RESULT1[60]), 
        .SI(MESSAGE1[60]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[140]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_141_ ( .D(RESULT1[61]), 
        .SI(MESSAGE1[61]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[141]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_142_ ( .D(RESULT1[62]), 
        .SI(MESSAGE1[62]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[142]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_143_ ( .D(RESULT1[63]), 
        .SI(MESSAGE1[63]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[143]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_144_ ( .D(RESULT1[48]), 
        .SI(MESSAGE1[48]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[144]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_145_ ( .D(RESULT1[49]), 
        .SI(MESSAGE1[49]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[145]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_146_ ( .D(RESULT1[50]), 
        .SI(MESSAGE1[50]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[146]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_147_ ( .D(RESULT1[51]), 
        .SI(MESSAGE1[51]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[147]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_148_ ( .D(RESULT1[52]), 
        .SI(MESSAGE1[52]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[148]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_149_ ( .D(RESULT1[53]), 
        .SI(MESSAGE1[53]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[149]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_150_ ( .D(RESULT1[54]), 
        .SI(MESSAGE1[54]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[150]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_151_ ( .D(RESULT1[55]), 
        .SI(MESSAGE1[55]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[151]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_152_ ( .D(RESULT1[40]), 
        .SI(MESSAGE1[40]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[152]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_153_ ( .D(RESULT1[41]), 
        .SI(MESSAGE1[41]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[153]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_154_ ( .D(RESULT1[42]), 
        .SI(MESSAGE1[42]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[154]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_155_ ( .D(RESULT1[43]), 
        .SI(MESSAGE1[43]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[155]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_156_ ( .D(RESULT1[44]), 
        .SI(MESSAGE1[44]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[156]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_157_ ( .D(RESULT1[45]), 
        .SI(MESSAGE1[45]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[157]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_158_ ( .D(RESULT1[46]), 
        .SI(MESSAGE1[46]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[158]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_159_ ( .D(RESULT1[47]), 
        .SI(MESSAGE1[47]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[159]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_160_ ( .D(RESULT1[32]), 
        .SI(MESSAGE1[32]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[160]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_161_ ( .D(RESULT1[33]), 
        .SI(MESSAGE1[33]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[161]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_162_ ( .D(RESULT1[34]), 
        .SI(MESSAGE1[34]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[162]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_163_ ( .D(RESULT1[35]), 
        .SI(MESSAGE1[35]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[163]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_164_ ( .D(RESULT1[36]), 
        .SI(MESSAGE1[36]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[164]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_165_ ( .D(RESULT1[37]), 
        .SI(MESSAGE1[37]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[165]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_166_ ( .D(RESULT1[38]), 
        .SI(MESSAGE1[38]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[166]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_167_ ( .D(RESULT1[39]), 
        .SI(MESSAGE1[39]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[167]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_168_ ( .D(RESULT1[24]), 
        .SI(MESSAGE1[24]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[168]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_169_ ( .D(RESULT1[25]), 
        .SI(MESSAGE1[25]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[169]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_170_ ( .D(RESULT1[26]), 
        .SI(MESSAGE1[26]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[170]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_171_ ( .D(RESULT1[27]), 
        .SI(MESSAGE1[27]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[171]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_172_ ( .D(RESULT1[28]), 
        .SI(MESSAGE1[28]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[172]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_173_ ( .D(RESULT1[29]), 
        .SI(MESSAGE1[29]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[173]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_174_ ( .D(RESULT1[30]), 
        .SI(MESSAGE1[30]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[174]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_175_ ( .D(RESULT1[31]), 
        .SI(MESSAGE1[31]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[175]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_176_ ( .D(RESULT1[16]), 
        .SI(MESSAGE1[16]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[176]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_177_ ( .D(RESULT1[17]), 
        .SI(MESSAGE1[17]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[177]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_178_ ( .D(RESULT1[18]), 
        .SI(MESSAGE1[18]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[178]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_179_ ( .D(RESULT1[19]), 
        .SI(MESSAGE1[19]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[179]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_180_ ( .D(RESULT1[20]), 
        .SI(MESSAGE1[20]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[180]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_181_ ( .D(RESULT1[21]), 
        .SI(MESSAGE1[21]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[181]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_182_ ( .D(RESULT1[22]), 
        .SI(MESSAGE1[22]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[182]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_183_ ( .D(RESULT1[23]), 
        .SI(MESSAGE1[23]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[183]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_184_ ( .D(RESULT1[8]), 
        .SI(MESSAGE1[8]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[184]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_185_ ( .D(RESULT1[9]), 
        .SI(MESSAGE1[9]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[185]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_186_ ( .D(RESULT1[10]), 
        .SI(MESSAGE1[10]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[186]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_187_ ( .D(RESULT1[11]), 
        .SI(MESSAGE1[11]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[187]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_188_ ( .D(RESULT1[12]), 
        .SI(MESSAGE1[12]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[188]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_189_ ( .D(RESULT1[13]), 
        .SI(MESSAGE1[13]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[189]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_190_ ( .D(RESULT1[14]), 
        .SI(MESSAGE1[14]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[190]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_191_ ( .D(RESULT1[15]), 
        .SI(MESSAGE1[15]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[191]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_192_ ( .D(RESULT1[0]), 
        .SI(MESSAGE1[0]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[192]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_193_ ( .D(RESULT1[1]), 
        .SI(MESSAGE1[1]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[193]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_194_ ( .D(RESULT1[2]), 
        .SI(MESSAGE1[2]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[194]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_195_ ( .D(RESULT1[3]), 
        .SI(MESSAGE1[3]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[195]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_196_ ( .D(RESULT1[4]), 
        .SI(MESSAGE1[4]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[196]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_197_ ( .D(RESULT1[5]), 
        .SI(MESSAGE1[5]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[197]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_198_ ( .D(RESULT1[6]), 
        .SI(MESSAGE1[6]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[198]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg1_s_current_state_reg_199_ ( .D(RESULT1[7]), 
        .SI(MESSAGE1[7]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE1[199]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_0_ ( .D(RESULT2[192]), 
        .SI(MESSAGE2[192]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[0]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_1_ ( .D(RESULT2[193]), 
        .SI(MESSAGE2[193]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[1]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_2_ ( .D(RESULT2[194]), 
        .SI(MESSAGE2[194]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[2]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_3_ ( .D(RESULT2[195]), 
        .SI(MESSAGE2[195]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[3]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_4_ ( .D(RESULT2[196]), 
        .SI(MESSAGE2[196]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[4]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_5_ ( .D(RESULT2[197]), 
        .SI(MESSAGE2[197]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[5]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_6_ ( .D(RESULT2[198]), 
        .SI(MESSAGE2[198]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[6]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_7_ ( .D(RESULT2[199]), 
        .SI(MESSAGE2[199]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[7]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_8_ ( .D(RESULT2[184]), 
        .SI(MESSAGE2[184]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[8]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_9_ ( .D(RESULT2[185]), 
        .SI(MESSAGE2[185]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[9]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_10_ ( .D(RESULT2[186]), 
        .SI(MESSAGE2[186]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[10]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_11_ ( .D(RESULT2[187]), 
        .SI(MESSAGE2[187]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[11]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_12_ ( .D(RESULT2[188]), 
        .SI(MESSAGE2[188]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[12]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_13_ ( .D(RESULT2[189]), 
        .SI(MESSAGE2[189]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[13]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_14_ ( .D(RESULT2[190]), 
        .SI(MESSAGE2[190]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[14]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_15_ ( .D(RESULT2[191]), 
        .SI(MESSAGE2[191]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[15]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_16_ ( .D(RESULT2[176]), 
        .SI(MESSAGE2[176]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[16]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_17_ ( .D(RESULT2[177]), 
        .SI(MESSAGE2[177]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[17]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_18_ ( .D(RESULT2[178]), 
        .SI(MESSAGE2[178]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[18]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_19_ ( .D(RESULT2[179]), 
        .SI(MESSAGE2[179]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[19]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_20_ ( .D(RESULT2[180]), 
        .SI(MESSAGE2[180]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[20]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_21_ ( .D(RESULT2[181]), 
        .SI(MESSAGE2[181]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[21]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_22_ ( .D(RESULT2[182]), 
        .SI(MESSAGE2[182]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[22]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_23_ ( .D(RESULT2[183]), 
        .SI(MESSAGE2[183]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[23]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_24_ ( .D(RESULT2[168]), 
        .SI(MESSAGE2[168]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[24]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_25_ ( .D(RESULT2[169]), 
        .SI(MESSAGE2[169]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[25]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_26_ ( .D(RESULT2[170]), 
        .SI(MESSAGE2[170]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[26]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_27_ ( .D(RESULT2[171]), 
        .SI(MESSAGE2[171]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[27]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_28_ ( .D(RESULT2[172]), 
        .SI(MESSAGE2[172]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[28]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_29_ ( .D(RESULT2[173]), 
        .SI(MESSAGE2[173]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[29]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_30_ ( .D(RESULT2[174]), 
        .SI(MESSAGE2[174]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[30]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_31_ ( .D(RESULT2[175]), 
        .SI(MESSAGE2[175]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[31]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_32_ ( .D(RESULT2[160]), 
        .SI(MESSAGE2[160]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[32]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_33_ ( .D(RESULT2[161]), 
        .SI(MESSAGE2[161]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[33]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_34_ ( .D(RESULT2[162]), 
        .SI(MESSAGE2[162]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[34]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_35_ ( .D(RESULT2[163]), 
        .SI(MESSAGE2[163]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[35]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_36_ ( .D(RESULT2[164]), 
        .SI(MESSAGE2[164]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[36]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_37_ ( .D(RESULT2[165]), 
        .SI(MESSAGE2[165]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[37]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_38_ ( .D(RESULT2[166]), 
        .SI(MESSAGE2[166]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[38]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_39_ ( .D(RESULT2[167]), 
        .SI(MESSAGE2[167]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[39]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_40_ ( .D(RESULT2[152]), 
        .SI(MESSAGE2[152]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[40]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_41_ ( .D(RESULT2[153]), 
        .SI(MESSAGE2[153]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[41]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_42_ ( .D(RESULT2[154]), 
        .SI(MESSAGE2[154]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[42]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_43_ ( .D(RESULT2[155]), 
        .SI(MESSAGE2[155]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[43]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_44_ ( .D(RESULT2[156]), 
        .SI(MESSAGE2[156]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[44]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_45_ ( .D(RESULT2[157]), 
        .SI(MESSAGE2[157]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[45]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_46_ ( .D(RESULT2[158]), 
        .SI(MESSAGE2[158]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[46]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_47_ ( .D(RESULT2[159]), 
        .SI(MESSAGE2[159]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[47]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_48_ ( .D(RESULT2[144]), 
        .SI(MESSAGE2[144]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[48]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_49_ ( .D(RESULT2[145]), 
        .SI(MESSAGE2[145]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[49]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_50_ ( .D(RESULT2[146]), 
        .SI(MESSAGE2[146]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[50]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_51_ ( .D(RESULT2[147]), 
        .SI(MESSAGE2[147]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[51]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_52_ ( .D(RESULT2[148]), 
        .SI(MESSAGE2[148]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[52]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_53_ ( .D(RESULT2[149]), 
        .SI(MESSAGE2[149]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[53]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_54_ ( .D(RESULT2[150]), 
        .SI(MESSAGE2[150]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[54]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_55_ ( .D(RESULT2[151]), 
        .SI(MESSAGE2[151]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[55]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_56_ ( .D(RESULT2[136]), 
        .SI(MESSAGE2[136]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[56]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_57_ ( .D(RESULT2[137]), 
        .SI(MESSAGE2[137]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[57]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_58_ ( .D(RESULT2[138]), 
        .SI(MESSAGE2[138]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[58]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_59_ ( .D(RESULT2[139]), 
        .SI(MESSAGE2[139]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[59]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_60_ ( .D(RESULT2[140]), 
        .SI(MESSAGE2[140]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[60]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_61_ ( .D(RESULT2[141]), 
        .SI(MESSAGE2[141]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[61]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_62_ ( .D(RESULT2[142]), 
        .SI(MESSAGE2[142]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[62]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_63_ ( .D(RESULT2[143]), 
        .SI(MESSAGE2[143]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[63]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_64_ ( .D(RESULT2[128]), 
        .SI(MESSAGE2[128]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[64]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_65_ ( .D(RESULT2[129]), 
        .SI(MESSAGE2[129]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[65]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_66_ ( .D(RESULT2[130]), 
        .SI(MESSAGE2[130]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[66]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_67_ ( .D(RESULT2[131]), 
        .SI(MESSAGE2[131]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[67]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_68_ ( .D(RESULT2[132]), 
        .SI(MESSAGE2[132]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[68]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_69_ ( .D(RESULT2[133]), 
        .SI(MESSAGE2[133]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[69]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_70_ ( .D(RESULT2[134]), 
        .SI(MESSAGE2[134]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[70]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_71_ ( .D(RESULT2[135]), 
        .SI(MESSAGE2[135]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[71]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_72_ ( .D(RESULT2[120]), 
        .SI(MESSAGE2[120]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[72]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_73_ ( .D(RESULT2[121]), 
        .SI(MESSAGE2[121]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[73]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_74_ ( .D(RESULT2[122]), 
        .SI(MESSAGE2[122]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[74]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_75_ ( .D(RESULT2[123]), 
        .SI(MESSAGE2[123]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[75]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_76_ ( .D(RESULT2[124]), 
        .SI(MESSAGE2[124]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[76]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_77_ ( .D(RESULT2[125]), 
        .SI(MESSAGE2[125]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[77]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_78_ ( .D(RESULT2[126]), 
        .SI(MESSAGE2[126]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[78]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_79_ ( .D(RESULT2[127]), 
        .SI(MESSAGE2[127]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[79]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_80_ ( .D(RESULT2[112]), 
        .SI(MESSAGE2[112]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[80]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_81_ ( .D(RESULT2[113]), 
        .SI(MESSAGE2[113]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[81]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_82_ ( .D(RESULT2[114]), 
        .SI(MESSAGE2[114]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[82]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_83_ ( .D(RESULT2[115]), 
        .SI(MESSAGE2[115]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[83]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_84_ ( .D(RESULT2[116]), 
        .SI(MESSAGE2[116]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[84]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_85_ ( .D(RESULT2[117]), 
        .SI(MESSAGE2[117]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[85]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_86_ ( .D(RESULT2[118]), 
        .SI(MESSAGE2[118]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[86]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_87_ ( .D(RESULT2[119]), 
        .SI(MESSAGE2[119]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[87]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_88_ ( .D(RESULT2[104]), 
        .SI(MESSAGE2[104]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[88]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_89_ ( .D(RESULT2[105]), 
        .SI(MESSAGE2[105]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[89]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_90_ ( .D(RESULT2[106]), 
        .SI(MESSAGE2[106]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[90]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_91_ ( .D(RESULT2[107]), 
        .SI(MESSAGE2[107]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[91]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_92_ ( .D(RESULT2[108]), 
        .SI(MESSAGE2[108]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[92]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_93_ ( .D(RESULT2[109]), 
        .SI(MESSAGE2[109]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[93]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_94_ ( .D(RESULT2[110]), 
        .SI(MESSAGE2[110]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[94]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_95_ ( .D(RESULT2[111]), 
        .SI(MESSAGE2[111]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[95]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_96_ ( .D(RESULT2[96]), 
        .SI(MESSAGE2[96]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[96]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_97_ ( .D(RESULT2[97]), 
        .SI(MESSAGE2[97]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[97]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_98_ ( .D(RESULT2[98]), 
        .SI(MESSAGE2[98]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[98]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_99_ ( .D(RESULT2[99]), 
        .SI(MESSAGE2[99]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[99]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_100_ ( .D(RESULT2[100]), 
        .SI(MESSAGE2[100]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[100]), .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_101_ ( .D(RESULT2[101]), 
        .SI(MESSAGE2[101]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[101]), .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_102_ ( .D(RESULT2[102]), 
        .SI(MESSAGE2[102]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[102]), .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_103_ ( .D(RESULT2[103]), 
        .SI(MESSAGE2[103]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[103]), .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_104_ ( .D(RESULT2[88]), 
        .SI(MESSAGE2[88]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[104]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_105_ ( .D(RESULT2[89]), 
        .SI(MESSAGE2[89]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[105]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_106_ ( .D(RESULT2[90]), 
        .SI(MESSAGE2[90]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[106]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_107_ ( .D(RESULT2[91]), 
        .SI(MESSAGE2[91]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[107]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_108_ ( .D(RESULT2[92]), 
        .SI(MESSAGE2[92]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[108]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_109_ ( .D(RESULT2[93]), 
        .SI(MESSAGE2[93]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[109]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_110_ ( .D(RESULT2[94]), 
        .SI(MESSAGE2[94]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[110]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_111_ ( .D(RESULT2[95]), 
        .SI(MESSAGE2[95]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[111]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_112_ ( .D(RESULT2[80]), 
        .SI(MESSAGE2[80]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[112]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_113_ ( .D(RESULT2[81]), 
        .SI(MESSAGE2[81]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[113]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_114_ ( .D(RESULT2[82]), 
        .SI(MESSAGE2[82]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[114]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_115_ ( .D(RESULT2[83]), 
        .SI(MESSAGE2[83]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[115]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_116_ ( .D(RESULT2[84]), 
        .SI(MESSAGE2[84]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[116]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_117_ ( .D(RESULT2[85]), 
        .SI(MESSAGE2[85]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[117]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_118_ ( .D(RESULT2[86]), 
        .SI(MESSAGE2[86]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[118]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_119_ ( .D(RESULT2[87]), 
        .SI(MESSAGE2[87]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[119]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_120_ ( .D(RESULT2[72]), 
        .SI(MESSAGE2[72]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[120]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_121_ ( .D(RESULT2[73]), 
        .SI(MESSAGE2[73]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[121]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_122_ ( .D(RESULT2[74]), 
        .SI(MESSAGE2[74]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[122]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_123_ ( .D(RESULT2[75]), 
        .SI(MESSAGE2[75]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[123]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_124_ ( .D(RESULT2[76]), 
        .SI(MESSAGE2[76]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[124]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_125_ ( .D(RESULT2[77]), 
        .SI(MESSAGE2[77]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[125]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_126_ ( .D(RESULT2[78]), 
        .SI(MESSAGE2[78]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[126]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_127_ ( .D(RESULT2[79]), 
        .SI(MESSAGE2[79]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[127]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_128_ ( .D(RESULT2[64]), 
        .SI(MESSAGE2[64]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[128]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_129_ ( .D(RESULT2[65]), 
        .SI(MESSAGE2[65]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[129]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_130_ ( .D(RESULT2[66]), 
        .SI(MESSAGE2[66]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[130]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_131_ ( .D(RESULT2[67]), 
        .SI(MESSAGE2[67]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[131]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_132_ ( .D(RESULT2[68]), 
        .SI(MESSAGE2[68]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[132]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_133_ ( .D(RESULT2[69]), 
        .SI(MESSAGE2[69]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[133]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_134_ ( .D(RESULT2[70]), 
        .SI(MESSAGE2[70]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[134]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_135_ ( .D(RESULT2[71]), 
        .SI(MESSAGE2[71]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[135]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_136_ ( .D(RESULT2[56]), 
        .SI(MESSAGE2[56]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[136]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_137_ ( .D(RESULT2[57]), 
        .SI(MESSAGE2[57]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[137]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_138_ ( .D(RESULT2[58]), 
        .SI(MESSAGE2[58]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[138]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_139_ ( .D(RESULT2[59]), 
        .SI(MESSAGE2[59]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[139]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_140_ ( .D(RESULT2[60]), 
        .SI(MESSAGE2[60]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[140]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_141_ ( .D(RESULT2[61]), 
        .SI(MESSAGE2[61]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[141]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_142_ ( .D(RESULT2[62]), 
        .SI(MESSAGE2[62]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[142]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_143_ ( .D(RESULT2[63]), 
        .SI(MESSAGE2[63]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[143]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_144_ ( .D(RESULT2[48]), 
        .SI(MESSAGE2[48]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[144]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_145_ ( .D(RESULT2[49]), 
        .SI(MESSAGE2[49]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[145]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_146_ ( .D(RESULT2[50]), 
        .SI(MESSAGE2[50]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[146]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_147_ ( .D(RESULT2[51]), 
        .SI(MESSAGE2[51]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[147]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_148_ ( .D(RESULT2[52]), 
        .SI(MESSAGE2[52]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[148]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_149_ ( .D(RESULT2[53]), 
        .SI(MESSAGE2[53]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[149]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_150_ ( .D(RESULT2[54]), 
        .SI(MESSAGE2[54]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[150]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_151_ ( .D(RESULT2[55]), 
        .SI(MESSAGE2[55]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[151]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_152_ ( .D(RESULT2[40]), 
        .SI(MESSAGE2[40]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[152]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_153_ ( .D(RESULT2[41]), 
        .SI(MESSAGE2[41]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[153]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_154_ ( .D(RESULT2[42]), 
        .SI(MESSAGE2[42]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[154]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_155_ ( .D(RESULT2[43]), 
        .SI(MESSAGE2[43]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[155]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_156_ ( .D(RESULT2[44]), 
        .SI(MESSAGE2[44]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[156]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_157_ ( .D(RESULT2[45]), 
        .SI(MESSAGE2[45]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[157]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_158_ ( .D(RESULT2[46]), 
        .SI(MESSAGE2[46]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[158]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_159_ ( .D(RESULT2[47]), 
        .SI(MESSAGE2[47]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[159]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_160_ ( .D(RESULT2[32]), 
        .SI(MESSAGE2[32]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[160]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_161_ ( .D(RESULT2[33]), 
        .SI(MESSAGE2[33]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[161]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_162_ ( .D(RESULT2[34]), 
        .SI(MESSAGE2[34]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[162]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_163_ ( .D(RESULT2[35]), 
        .SI(MESSAGE2[35]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[163]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_164_ ( .D(RESULT2[36]), 
        .SI(MESSAGE2[36]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[164]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_165_ ( .D(RESULT2[37]), 
        .SI(MESSAGE2[37]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[165]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_166_ ( .D(RESULT2[38]), 
        .SI(MESSAGE2[38]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[166]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_167_ ( .D(RESULT2[39]), 
        .SI(MESSAGE2[39]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[167]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_168_ ( .D(RESULT2[24]), 
        .SI(MESSAGE2[24]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[168]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_169_ ( .D(RESULT2[25]), 
        .SI(MESSAGE2[25]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[169]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_170_ ( .D(RESULT2[26]), 
        .SI(MESSAGE2[26]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[170]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_171_ ( .D(RESULT2[27]), 
        .SI(MESSAGE2[27]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[171]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_172_ ( .D(RESULT2[28]), 
        .SI(MESSAGE2[28]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[172]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_173_ ( .D(RESULT2[29]), 
        .SI(MESSAGE2[29]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[173]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_174_ ( .D(RESULT2[30]), 
        .SI(MESSAGE2[30]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[174]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_175_ ( .D(RESULT2[31]), 
        .SI(MESSAGE2[31]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[175]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_176_ ( .D(RESULT2[16]), 
        .SI(MESSAGE2[16]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[176]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_177_ ( .D(RESULT2[17]), 
        .SI(MESSAGE2[17]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[177]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_178_ ( .D(RESULT2[18]), 
        .SI(MESSAGE2[18]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[178]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_179_ ( .D(RESULT2[19]), 
        .SI(MESSAGE2[19]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[179]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_180_ ( .D(RESULT2[20]), 
        .SI(MESSAGE2[20]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[180]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_181_ ( .D(RESULT2[21]), 
        .SI(MESSAGE2[21]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[181]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_182_ ( .D(RESULT2[22]), 
        .SI(MESSAGE2[22]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[182]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_183_ ( .D(RESULT2[23]), 
        .SI(MESSAGE2[23]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[183]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_184_ ( .D(RESULT2[8]), 
        .SI(MESSAGE2[8]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[184]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_185_ ( .D(RESULT2[9]), 
        .SI(MESSAGE2[9]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[185]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_186_ ( .D(RESULT2[10]), 
        .SI(MESSAGE2[10]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[186]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_187_ ( .D(RESULT2[11]), 
        .SI(MESSAGE2[11]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[187]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_188_ ( .D(RESULT2[12]), 
        .SI(MESSAGE2[12]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[188]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_189_ ( .D(RESULT2[13]), 
        .SI(MESSAGE2[13]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[189]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_190_ ( .D(RESULT2[14]), 
        .SI(MESSAGE2[14]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[190]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_191_ ( .D(RESULT2[15]), 
        .SI(MESSAGE2[15]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[191]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_192_ ( .D(RESULT2[0]), 
        .SI(MESSAGE2[0]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[192]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_193_ ( .D(RESULT2[1]), 
        .SI(MESSAGE2[1]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[193]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_194_ ( .D(RESULT2[2]), 
        .SI(MESSAGE2[2]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[194]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_195_ ( .D(RESULT2[3]), 
        .SI(MESSAGE2[3]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[195]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_196_ ( .D(RESULT2[4]), 
        .SI(MESSAGE2[4]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[196]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_197_ ( .D(RESULT2[5]), 
        .SI(MESSAGE2[5]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[197]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_198_ ( .D(RESULT2[6]), 
        .SI(MESSAGE2[6]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[198]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg2_s_current_state_reg_199_ ( .D(RESULT2[7]), 
        .SI(MESSAGE2[7]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE2[199]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_0_ ( .D(RESULT3[192]), 
        .SI(MESSAGE3[192]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[0]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_1_ ( .D(RESULT3[193]), 
        .SI(MESSAGE3[193]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[1]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_2_ ( .D(RESULT3[194]), 
        .SI(MESSAGE3[194]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[2]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_3_ ( .D(RESULT3[195]), 
        .SI(MESSAGE3[195]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[3]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_4_ ( .D(RESULT3[196]), 
        .SI(MESSAGE3[196]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[4]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_5_ ( .D(RESULT3[197]), 
        .SI(MESSAGE3[197]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[5]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_6_ ( .D(RESULT3[198]), 
        .SI(MESSAGE3[198]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[6]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_7_ ( .D(RESULT3[199]), 
        .SI(MESSAGE3[199]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[7]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_8_ ( .D(RESULT3[184]), 
        .SI(MESSAGE3[184]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[8]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_9_ ( .D(RESULT3[185]), 
        .SI(MESSAGE3[185]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[9]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_10_ ( .D(RESULT3[186]), 
        .SI(MESSAGE3[186]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[10]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_11_ ( .D(RESULT3[187]), 
        .SI(MESSAGE3[187]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[11]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_12_ ( .D(RESULT3[188]), 
        .SI(MESSAGE3[188]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[12]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_13_ ( .D(RESULT3[189]), 
        .SI(MESSAGE3[189]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[13]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_14_ ( .D(RESULT3[190]), 
        .SI(MESSAGE3[190]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[14]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_15_ ( .D(RESULT3[191]), 
        .SI(MESSAGE3[191]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[15]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_16_ ( .D(RESULT3[176]), 
        .SI(MESSAGE3[176]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[16]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_17_ ( .D(RESULT3[177]), 
        .SI(MESSAGE3[177]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[17]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_18_ ( .D(RESULT3[178]), 
        .SI(MESSAGE3[178]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[18]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_19_ ( .D(RESULT3[179]), 
        .SI(MESSAGE3[179]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[19]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_20_ ( .D(RESULT3[180]), 
        .SI(MESSAGE3[180]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[20]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_21_ ( .D(RESULT3[181]), 
        .SI(MESSAGE3[181]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[21]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_22_ ( .D(RESULT3[182]), 
        .SI(MESSAGE3[182]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[22]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_23_ ( .D(RESULT3[183]), 
        .SI(MESSAGE3[183]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[23]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_24_ ( .D(RESULT3[168]), 
        .SI(MESSAGE3[168]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[24]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_25_ ( .D(RESULT3[169]), 
        .SI(MESSAGE3[169]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[25]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_26_ ( .D(RESULT3[170]), 
        .SI(MESSAGE3[170]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[26]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_27_ ( .D(RESULT3[171]), 
        .SI(MESSAGE3[171]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[27]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_28_ ( .D(RESULT3[172]), 
        .SI(MESSAGE3[172]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[28]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_29_ ( .D(RESULT3[173]), 
        .SI(MESSAGE3[173]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[29]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_30_ ( .D(RESULT3[174]), 
        .SI(MESSAGE3[174]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[30]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_31_ ( .D(RESULT3[175]), 
        .SI(MESSAGE3[175]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[31]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_32_ ( .D(RESULT3[160]), 
        .SI(MESSAGE3[160]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[32]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_33_ ( .D(RESULT3[161]), 
        .SI(MESSAGE3[161]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[33]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_34_ ( .D(RESULT3[162]), 
        .SI(MESSAGE3[162]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[34]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_35_ ( .D(RESULT3[163]), 
        .SI(MESSAGE3[163]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[35]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_36_ ( .D(RESULT3[164]), 
        .SI(MESSAGE3[164]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[36]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_37_ ( .D(RESULT3[165]), 
        .SI(MESSAGE3[165]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[37]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_38_ ( .D(RESULT3[166]), 
        .SI(MESSAGE3[166]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[38]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_39_ ( .D(RESULT3[167]), 
        .SI(MESSAGE3[167]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[39]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_40_ ( .D(RESULT3[152]), 
        .SI(MESSAGE3[152]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[40]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_41_ ( .D(RESULT3[153]), 
        .SI(MESSAGE3[153]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[41]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_42_ ( .D(RESULT3[154]), 
        .SI(MESSAGE3[154]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[42]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_43_ ( .D(RESULT3[155]), 
        .SI(MESSAGE3[155]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[43]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_44_ ( .D(RESULT3[156]), 
        .SI(MESSAGE3[156]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[44]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_45_ ( .D(RESULT3[157]), 
        .SI(MESSAGE3[157]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[45]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_46_ ( .D(RESULT3[158]), 
        .SI(MESSAGE3[158]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[46]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_47_ ( .D(RESULT3[159]), 
        .SI(MESSAGE3[159]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[47]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_48_ ( .D(RESULT3[144]), 
        .SI(MESSAGE3[144]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[48]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_49_ ( .D(RESULT3[145]), 
        .SI(MESSAGE3[145]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[49]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_50_ ( .D(RESULT3[146]), 
        .SI(MESSAGE3[146]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[50]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_51_ ( .D(RESULT3[147]), 
        .SI(MESSAGE3[147]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[51]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_52_ ( .D(RESULT3[148]), 
        .SI(MESSAGE3[148]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[52]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_53_ ( .D(RESULT3[149]), 
        .SI(MESSAGE3[149]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[53]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_54_ ( .D(RESULT3[150]), 
        .SI(MESSAGE3[150]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[54]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_55_ ( .D(RESULT3[151]), 
        .SI(MESSAGE3[151]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[55]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_56_ ( .D(RESULT3[136]), 
        .SI(MESSAGE3[136]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[56]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_57_ ( .D(RESULT3[137]), 
        .SI(MESSAGE3[137]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[57]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_58_ ( .D(RESULT3[138]), 
        .SI(MESSAGE3[138]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[58]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_59_ ( .D(RESULT3[139]), 
        .SI(MESSAGE3[139]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[59]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_60_ ( .D(RESULT3[140]), 
        .SI(MESSAGE3[140]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[60]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_61_ ( .D(RESULT3[141]), 
        .SI(MESSAGE3[141]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[61]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_62_ ( .D(RESULT3[142]), 
        .SI(MESSAGE3[142]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[62]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_63_ ( .D(RESULT3[143]), 
        .SI(MESSAGE3[143]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[63]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_64_ ( .D(RESULT3[128]), 
        .SI(MESSAGE3[128]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[64]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_65_ ( .D(RESULT3[129]), 
        .SI(MESSAGE3[129]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[65]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_66_ ( .D(RESULT3[130]), 
        .SI(MESSAGE3[130]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[66]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_67_ ( .D(RESULT3[131]), 
        .SI(MESSAGE3[131]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[67]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_68_ ( .D(RESULT3[132]), 
        .SI(MESSAGE3[132]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[68]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_69_ ( .D(RESULT3[133]), 
        .SI(MESSAGE3[133]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[69]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_70_ ( .D(RESULT3[134]), 
        .SI(MESSAGE3[134]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[70]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_71_ ( .D(RESULT3[135]), 
        .SI(MESSAGE3[135]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[71]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_72_ ( .D(RESULT3[120]), 
        .SI(MESSAGE3[120]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[72]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_73_ ( .D(RESULT3[121]), 
        .SI(MESSAGE3[121]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[73]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_74_ ( .D(RESULT3[122]), 
        .SI(MESSAGE3[122]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[74]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_75_ ( .D(RESULT3[123]), 
        .SI(MESSAGE3[123]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[75]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_76_ ( .D(RESULT3[124]), 
        .SI(MESSAGE3[124]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[76]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_77_ ( .D(RESULT3[125]), 
        .SI(MESSAGE3[125]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[77]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_78_ ( .D(RESULT3[126]), 
        .SI(MESSAGE3[126]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[78]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_79_ ( .D(RESULT3[127]), 
        .SI(MESSAGE3[127]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[79]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_80_ ( .D(RESULT3[112]), 
        .SI(MESSAGE3[112]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[80]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_81_ ( .D(RESULT3[113]), 
        .SI(MESSAGE3[113]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[81]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_82_ ( .D(RESULT3[114]), 
        .SI(MESSAGE3[114]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[82]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_83_ ( .D(RESULT3[115]), 
        .SI(MESSAGE3[115]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[83]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_84_ ( .D(RESULT3[116]), 
        .SI(MESSAGE3[116]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[84]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_85_ ( .D(RESULT3[117]), 
        .SI(MESSAGE3[117]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[85]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_86_ ( .D(RESULT3[118]), 
        .SI(MESSAGE3[118]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[86]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_87_ ( .D(RESULT3[119]), 
        .SI(MESSAGE3[119]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[87]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_88_ ( .D(RESULT3[104]), 
        .SI(MESSAGE3[104]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[88]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_89_ ( .D(RESULT3[105]), 
        .SI(MESSAGE3[105]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[89]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_90_ ( .D(RESULT3[106]), 
        .SI(MESSAGE3[106]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[90]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_91_ ( .D(RESULT3[107]), 
        .SI(MESSAGE3[107]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[91]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_92_ ( .D(RESULT3[108]), 
        .SI(MESSAGE3[108]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[92]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_93_ ( .D(RESULT3[109]), 
        .SI(MESSAGE3[109]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[93]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_94_ ( .D(RESULT3[110]), 
        .SI(MESSAGE3[110]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[94]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_95_ ( .D(RESULT3[111]), 
        .SI(MESSAGE3[111]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[95]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_96_ ( .D(RESULT3[96]), 
        .SI(MESSAGE3[96]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[96]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_97_ ( .D(RESULT3[97]), 
        .SI(MESSAGE3[97]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[97]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_98_ ( .D(RESULT3[98]), 
        .SI(MESSAGE3[98]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[98]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_99_ ( .D(RESULT3[99]), 
        .SI(MESSAGE3[99]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[99]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_100_ ( .D(RESULT3[100]), 
        .SI(MESSAGE3[100]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[100]), .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_101_ ( .D(RESULT3[101]), 
        .SI(MESSAGE3[101]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[101]), .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_102_ ( .D(RESULT3[102]), 
        .SI(MESSAGE3[102]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[102]), .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_103_ ( .D(RESULT3[103]), 
        .SI(MESSAGE3[103]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[103]), .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_104_ ( .D(RESULT3[88]), 
        .SI(MESSAGE3[88]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[104]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_105_ ( .D(RESULT3[89]), 
        .SI(MESSAGE3[89]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[105]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_106_ ( .D(RESULT3[90]), 
        .SI(MESSAGE3[90]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[106]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_107_ ( .D(RESULT3[91]), 
        .SI(MESSAGE3[91]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[107]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_108_ ( .D(RESULT3[92]), 
        .SI(MESSAGE3[92]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[108]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_109_ ( .D(RESULT3[93]), 
        .SI(MESSAGE3[93]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[109]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_110_ ( .D(RESULT3[94]), 
        .SI(MESSAGE3[94]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[110]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_111_ ( .D(RESULT3[95]), 
        .SI(MESSAGE3[95]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[111]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_112_ ( .D(RESULT3[80]), 
        .SI(MESSAGE3[80]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[112]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_113_ ( .D(RESULT3[81]), 
        .SI(MESSAGE3[81]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[113]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_114_ ( .D(RESULT3[82]), 
        .SI(MESSAGE3[82]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[114]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_115_ ( .D(RESULT3[83]), 
        .SI(MESSAGE3[83]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[115]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_116_ ( .D(RESULT3[84]), 
        .SI(MESSAGE3[84]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[116]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_117_ ( .D(RESULT3[85]), 
        .SI(MESSAGE3[85]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[117]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_118_ ( .D(RESULT3[86]), 
        .SI(MESSAGE3[86]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[118]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_119_ ( .D(RESULT3[87]), 
        .SI(MESSAGE3[87]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[119]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_120_ ( .D(RESULT3[72]), 
        .SI(MESSAGE3[72]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[120]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_121_ ( .D(RESULT3[73]), 
        .SI(MESSAGE3[73]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[121]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_122_ ( .D(RESULT3[74]), 
        .SI(MESSAGE3[74]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[122]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_123_ ( .D(RESULT3[75]), 
        .SI(MESSAGE3[75]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[123]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_124_ ( .D(RESULT3[76]), 
        .SI(MESSAGE3[76]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[124]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_125_ ( .D(RESULT3[77]), 
        .SI(MESSAGE3[77]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[125]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_126_ ( .D(RESULT3[78]), 
        .SI(MESSAGE3[78]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[126]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_127_ ( .D(RESULT3[79]), 
        .SI(MESSAGE3[79]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[127]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_128_ ( .D(RESULT3[64]), 
        .SI(MESSAGE3[64]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[128]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_129_ ( .D(RESULT3[65]), 
        .SI(MESSAGE3[65]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[129]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_130_ ( .D(RESULT3[66]), 
        .SI(MESSAGE3[66]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[130]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_131_ ( .D(RESULT3[67]), 
        .SI(MESSAGE3[67]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[131]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_132_ ( .D(RESULT3[68]), 
        .SI(MESSAGE3[68]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[132]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_133_ ( .D(RESULT3[69]), 
        .SI(MESSAGE3[69]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[133]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_134_ ( .D(RESULT3[70]), 
        .SI(MESSAGE3[70]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[134]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_135_ ( .D(RESULT3[71]), 
        .SI(MESSAGE3[71]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[135]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_136_ ( .D(RESULT3[56]), 
        .SI(MESSAGE3[56]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[136]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_137_ ( .D(RESULT3[57]), 
        .SI(MESSAGE3[57]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[137]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_138_ ( .D(RESULT3[58]), 
        .SI(MESSAGE3[58]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[138]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_139_ ( .D(RESULT3[59]), 
        .SI(MESSAGE3[59]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[139]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_140_ ( .D(RESULT3[60]), 
        .SI(MESSAGE3[60]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[140]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_141_ ( .D(RESULT3[61]), 
        .SI(MESSAGE3[61]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[141]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_142_ ( .D(RESULT3[62]), 
        .SI(MESSAGE3[62]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[142]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_143_ ( .D(RESULT3[63]), 
        .SI(MESSAGE3[63]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[143]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_144_ ( .D(RESULT3[48]), 
        .SI(MESSAGE3[48]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[144]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_145_ ( .D(RESULT3[49]), 
        .SI(MESSAGE3[49]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[145]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_146_ ( .D(RESULT3[50]), 
        .SI(MESSAGE3[50]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[146]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_147_ ( .D(RESULT3[51]), 
        .SI(MESSAGE3[51]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[147]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_148_ ( .D(RESULT3[52]), 
        .SI(MESSAGE3[52]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[148]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_149_ ( .D(RESULT3[53]), 
        .SI(MESSAGE3[53]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[149]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_150_ ( .D(RESULT3[54]), 
        .SI(MESSAGE3[54]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[150]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_151_ ( .D(RESULT3[55]), 
        .SI(MESSAGE3[55]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[151]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_152_ ( .D(RESULT3[40]), 
        .SI(MESSAGE3[40]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[152]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_153_ ( .D(RESULT3[41]), 
        .SI(MESSAGE3[41]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[153]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_154_ ( .D(RESULT3[42]), 
        .SI(MESSAGE3[42]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[154]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_155_ ( .D(RESULT3[43]), 
        .SI(MESSAGE3[43]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[155]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_156_ ( .D(RESULT3[44]), 
        .SI(MESSAGE3[44]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[156]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_157_ ( .D(RESULT3[45]), 
        .SI(MESSAGE3[45]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[157]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_158_ ( .D(RESULT3[46]), 
        .SI(MESSAGE3[46]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[158]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_159_ ( .D(RESULT3[47]), 
        .SI(MESSAGE3[47]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[159]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_160_ ( .D(RESULT3[32]), 
        .SI(MESSAGE3[32]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[160]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_161_ ( .D(RESULT3[33]), 
        .SI(MESSAGE3[33]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[161]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_162_ ( .D(RESULT3[34]), 
        .SI(MESSAGE3[34]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[162]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_163_ ( .D(RESULT3[35]), 
        .SI(MESSAGE3[35]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[163]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_164_ ( .D(RESULT3[36]), 
        .SI(MESSAGE3[36]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[164]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_165_ ( .D(RESULT3[37]), 
        .SI(MESSAGE3[37]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[165]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_166_ ( .D(RESULT3[38]), 
        .SI(MESSAGE3[38]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[166]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_167_ ( .D(RESULT3[39]), 
        .SI(MESSAGE3[39]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[167]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_168_ ( .D(RESULT3[24]), 
        .SI(MESSAGE3[24]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[168]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_169_ ( .D(RESULT3[25]), 
        .SI(MESSAGE3[25]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[169]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_170_ ( .D(RESULT3[26]), 
        .SI(MESSAGE3[26]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[170]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_171_ ( .D(RESULT3[27]), 
        .SI(MESSAGE3[27]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[171]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_172_ ( .D(RESULT3[28]), 
        .SI(MESSAGE3[28]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[172]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_173_ ( .D(RESULT3[29]), 
        .SI(MESSAGE3[29]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[173]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_174_ ( .D(RESULT3[30]), 
        .SI(MESSAGE3[30]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[174]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_175_ ( .D(RESULT3[31]), 
        .SI(MESSAGE3[31]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[175]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_176_ ( .D(RESULT3[16]), 
        .SI(MESSAGE3[16]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[176]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_177_ ( .D(RESULT3[17]), 
        .SI(MESSAGE3[17]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[177]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_178_ ( .D(RESULT3[18]), 
        .SI(MESSAGE3[18]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[178]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_179_ ( .D(RESULT3[19]), 
        .SI(MESSAGE3[19]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[179]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_180_ ( .D(RESULT3[20]), 
        .SI(MESSAGE3[20]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[180]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_181_ ( .D(RESULT3[21]), 
        .SI(MESSAGE3[21]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[181]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_182_ ( .D(RESULT3[22]), 
        .SI(MESSAGE3[22]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[182]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_183_ ( .D(RESULT3[23]), 
        .SI(MESSAGE3[23]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[183]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_184_ ( .D(RESULT3[8]), 
        .SI(MESSAGE3[8]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[184]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_185_ ( .D(RESULT3[9]), 
        .SI(MESSAGE3[9]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[185]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_186_ ( .D(RESULT3[10]), 
        .SI(MESSAGE3[10]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[186]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_187_ ( .D(RESULT3[11]), 
        .SI(MESSAGE3[11]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[187]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_188_ ( .D(RESULT3[12]), 
        .SI(MESSAGE3[12]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[188]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_189_ ( .D(RESULT3[13]), 
        .SI(MESSAGE3[13]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[189]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_190_ ( .D(RESULT3[14]), 
        .SI(MESSAGE3[14]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[190]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_191_ ( .D(RESULT3[15]), 
        .SI(MESSAGE3[15]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[191]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_192_ ( .D(RESULT3[0]), 
        .SI(MESSAGE3[0]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[192]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_193_ ( .D(RESULT3[1]), 
        .SI(MESSAGE3[1]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[193]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_194_ ( .D(RESULT3[2]), 
        .SI(MESSAGE3[2]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[194]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_195_ ( .D(RESULT3[3]), 
        .SI(MESSAGE3[3]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[195]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_196_ ( .D(RESULT3[4]), 
        .SI(MESSAGE3[4]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[196]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_197_ ( .D(RESULT3[5]), 
        .SI(MESSAGE3[5]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[197]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_198_ ( .D(RESULT3[6]), 
        .SI(MESSAGE3[6]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[198]), 
        .QN() );
  SDFF_X1 RoundFunction_StateReg3_s_current_state_reg_199_ ( .D(RESULT3[7]), 
        .SI(MESSAGE3[7]), .SE(RESET), .CK(CLK), .Q(RoundFunction_STATE3[199]), 
        .QN() );
  XNOR2_X1 RoundFunction_T1_U400 ( .A(RoundFunction_STATE1[9]), .B(
        RoundFunction_T1_n600), .ZN(RoundFunction_TMP3_1[82]) );
  XNOR2_X1 RoundFunction_T1_U399 ( .A(RoundFunction_STATE1[99]), .B(
        RoundFunction_T1_n599), .ZN(RoundFunction_TMP3_1[22]) );
  XNOR2_X1 RoundFunction_T1_U398 ( .A(RoundFunction_STATE1[98]), .B(
        RoundFunction_T1_n598), .ZN(RoundFunction_TMP3_1[21]) );
  XNOR2_X1 RoundFunction_T1_U397 ( .A(RoundFunction_STATE1[97]), .B(
        RoundFunction_T1_n597), .ZN(RoundFunction_TMP3_1[20]) );
  XNOR2_X1 RoundFunction_T1_U396 ( .A(RoundFunction_STATE1[96]), .B(
        RoundFunction_T1_n596), .ZN(RoundFunction_TMP3_1[19]) );
  XNOR2_X1 RoundFunction_T1_U395 ( .A(RoundFunction_STATE1[95]), .B(
        RoundFunction_T1_n595), .ZN(RoundFunction_TMP3_1[137]) );
  XNOR2_X1 RoundFunction_T1_U394 ( .A(RoundFunction_STATE1[94]), .B(
        RoundFunction_T1_n594), .ZN(RoundFunction_TMP3_1[136]) );
  XNOR2_X1 RoundFunction_T1_U393 ( .A(RoundFunction_STATE1[93]), .B(
        RoundFunction_T1_n593), .ZN(RoundFunction_TMP3_1[143]) );
  XNOR2_X1 RoundFunction_T1_U392 ( .A(RoundFunction_STATE1[92]), .B(
        RoundFunction_T1_n592), .ZN(RoundFunction_TMP3_1[142]) );
  XNOR2_X1 RoundFunction_T1_U391 ( .A(RoundFunction_STATE1[91]), .B(
        RoundFunction_T1_n591), .ZN(RoundFunction_TMP3_1[141]) );
  XNOR2_X1 RoundFunction_T1_U390 ( .A(RoundFunction_STATE1[90]), .B(
        RoundFunction_T1_n590), .ZN(RoundFunction_TMP3_1[140]) );
  XNOR2_X1 RoundFunction_T1_U389 ( .A(RoundFunction_STATE1[8]), .B(
        RoundFunction_T1_n589), .ZN(RoundFunction_TMP3_1[81]) );
  XNOR2_X1 RoundFunction_T1_U388 ( .A(RoundFunction_STATE1[89]), .B(
        RoundFunction_T1_n600), .ZN(RoundFunction_TMP3_1[139]) );
  XNOR2_X1 RoundFunction_T1_U387 ( .A(RoundFunction_STATE1[88]), .B(
        RoundFunction_T1_n589), .ZN(RoundFunction_TMP3_1[138]) );
  XNOR2_X1 RoundFunction_T1_U386 ( .A(RoundFunction_STATE1[87]), .B(
        RoundFunction_T1_n588), .ZN(RoundFunction_TMP3_1[58]) );
  XNOR2_X1 RoundFunction_T1_U385 ( .A(RoundFunction_STATE1[86]), .B(
        RoundFunction_T1_n587), .ZN(RoundFunction_TMP3_1[57]) );
  XNOR2_X1 RoundFunction_T1_U384 ( .A(RoundFunction_STATE1[85]), .B(
        RoundFunction_T1_n586), .ZN(RoundFunction_TMP3_1[56]) );
  XNOR2_X1 RoundFunction_T1_U383 ( .A(RoundFunction_STATE1[84]), .B(
        RoundFunction_T1_n585), .ZN(RoundFunction_TMP3_1[63]) );
  XNOR2_X1 RoundFunction_T1_U382 ( .A(RoundFunction_STATE1[83]), .B(
        RoundFunction_T1_n584), .ZN(RoundFunction_TMP3_1[62]) );
  XNOR2_X1 RoundFunction_T1_U381 ( .A(RoundFunction_STATE1[82]), .B(
        RoundFunction_T1_n583), .ZN(RoundFunction_TMP3_1[61]) );
  XNOR2_X1 RoundFunction_T1_U380 ( .A(RoundFunction_STATE1[81]), .B(
        RoundFunction_T1_n582), .ZN(RoundFunction_TMP3_1[60]) );
  XNOR2_X1 RoundFunction_T1_U379 ( .A(RoundFunction_STATE1[80]), .B(
        RoundFunction_T1_n581), .ZN(RoundFunction_TMP3_1[59]) );
  XNOR2_X1 RoundFunction_T1_U378 ( .A(RoundFunction_STATE1[7]), .B(
        RoundFunction_T1_n588), .ZN(RoundFunction_TMP3_1[7]) );
  XNOR2_X1 RoundFunction_T1_U377 ( .A(RoundFunction_STATE1[79]), .B(
        RoundFunction_T1_n580), .ZN(RoundFunction_TMP3_1[51]) );
  XNOR2_X1 RoundFunction_T1_U376 ( .A(RoundFunction_STATE1[78]), .B(
        RoundFunction_T1_n579), .ZN(RoundFunction_TMP3_1[50]) );
  XNOR2_X1 RoundFunction_T1_U375 ( .A(RoundFunction_STATE1[77]), .B(
        RoundFunction_T1_n578), .ZN(RoundFunction_TMP3_1[49]) );
  XNOR2_X1 RoundFunction_T1_U374 ( .A(RoundFunction_STATE1[76]), .B(
        RoundFunction_T1_n577), .ZN(RoundFunction_TMP3_1[48]) );
  XNOR2_X1 RoundFunction_T1_U373 ( .A(RoundFunction_STATE1[75]), .B(
        RoundFunction_T1_n576), .ZN(RoundFunction_TMP3_1[55]) );
  XNOR2_X1 RoundFunction_T1_U372 ( .A(RoundFunction_STATE1[74]), .B(
        RoundFunction_T1_n575), .ZN(RoundFunction_TMP3_1[54]) );
  XNOR2_X1 RoundFunction_T1_U371 ( .A(RoundFunction_STATE1[73]), .B(
        RoundFunction_T1_n574), .ZN(RoundFunction_TMP3_1[53]) );
  XNOR2_X1 RoundFunction_T1_U370 ( .A(RoundFunction_STATE1[72]), .B(
        RoundFunction_T1_n573), .ZN(RoundFunction_TMP3_1[52]) );
  XNOR2_X1 RoundFunction_T1_U369 ( .A(RoundFunction_STATE1[71]), .B(
        RoundFunction_T1_n572), .ZN(RoundFunction_TMP3_1[174]) );
  XNOR2_X1 RoundFunction_T1_U368 ( .A(RoundFunction_STATE1[70]), .B(
        RoundFunction_T1_n571), .ZN(RoundFunction_TMP3_1[173]) );
  XNOR2_X1 RoundFunction_T1_U367 ( .A(RoundFunction_STATE1[6]), .B(
        RoundFunction_T1_n587), .ZN(RoundFunction_TMP3_1[6]) );
  XNOR2_X1 RoundFunction_T1_U366 ( .A(RoundFunction_STATE1[69]), .B(
        RoundFunction_T1_n570), .ZN(RoundFunction_TMP3_1[172]) );
  XNOR2_X1 RoundFunction_T1_U365 ( .A(RoundFunction_STATE1[68]), .B(
        RoundFunction_T1_n569), .ZN(RoundFunction_TMP3_1[171]) );
  XNOR2_X1 RoundFunction_T1_U364 ( .A(RoundFunction_STATE1[67]), .B(
        RoundFunction_T1_n568), .ZN(RoundFunction_TMP3_1[170]) );
  XNOR2_X1 RoundFunction_T1_U363 ( .A(RoundFunction_STATE1[66]), .B(
        RoundFunction_T1_n567), .ZN(RoundFunction_TMP3_1[169]) );
  XNOR2_X1 RoundFunction_T1_U362 ( .A(RoundFunction_STATE1[65]), .B(
        RoundFunction_T1_n566), .ZN(RoundFunction_TMP3_1[168]) );
  XNOR2_X1 RoundFunction_T1_U361 ( .A(RoundFunction_STATE1[64]), .B(
        RoundFunction_T1_n565), .ZN(RoundFunction_TMP3_1[175]) );
  XNOR2_X1 RoundFunction_T1_U360 ( .A(RoundFunction_STATE1[63]), .B(
        RoundFunction_T1_n564), .ZN(RoundFunction_TMP3_1[93]) );
  XNOR2_X1 RoundFunction_T1_U359 ( .A(RoundFunction_STATE1[62]), .B(
        RoundFunction_T1_n563), .ZN(RoundFunction_TMP3_1[92]) );
  XNOR2_X1 RoundFunction_T1_U358 ( .A(RoundFunction_STATE1[61]), .B(
        RoundFunction_T1_n562), .ZN(RoundFunction_TMP3_1[91]) );
  XNOR2_X1 RoundFunction_T1_U357 ( .A(RoundFunction_STATE1[60]), .B(
        RoundFunction_T1_n561), .ZN(RoundFunction_TMP3_1[90]) );
  XNOR2_X1 RoundFunction_T1_U356 ( .A(RoundFunction_STATE1[5]), .B(
        RoundFunction_T1_n586), .ZN(RoundFunction_TMP3_1[5]) );
  XNOR2_X1 RoundFunction_T1_U355 ( .A(RoundFunction_STATE1[59]), .B(
        RoundFunction_T1_n599), .ZN(RoundFunction_TMP3_1[89]) );
  XNOR2_X1 RoundFunction_T1_U354 ( .A(RoundFunction_STATE1[58]), .B(
        RoundFunction_T1_n598), .ZN(RoundFunction_TMP3_1[88]) );
  XNOR2_X1 RoundFunction_T1_U353 ( .A(RoundFunction_STATE1[57]), .B(
        RoundFunction_T1_n597), .ZN(RoundFunction_TMP3_1[95]) );
  XNOR2_X1 RoundFunction_T1_U352 ( .A(RoundFunction_STATE1[56]), .B(
        RoundFunction_T1_n596), .ZN(RoundFunction_TMP3_1[94]) );
  XNOR2_X1 RoundFunction_T1_U351 ( .A(RoundFunction_STATE1[55]), .B(
        RoundFunction_T1_n595), .ZN(RoundFunction_TMP3_1[11]) );
  XNOR2_X1 RoundFunction_T1_U350 ( .A(RoundFunction_STATE1[54]), .B(
        RoundFunction_T1_n594), .ZN(RoundFunction_TMP3_1[10]) );
  XNOR2_X1 RoundFunction_T1_U349 ( .A(RoundFunction_STATE1[53]), .B(
        RoundFunction_T1_n593), .ZN(RoundFunction_TMP3_1[9]) );
  XNOR2_X1 RoundFunction_T1_U348 ( .A(RoundFunction_STATE1[52]), .B(
        RoundFunction_T1_n592), .ZN(RoundFunction_TMP3_1[8]) );
  XNOR2_X1 RoundFunction_T1_U347 ( .A(RoundFunction_STATE1[51]), .B(
        RoundFunction_T1_n591), .ZN(RoundFunction_TMP3_1[15]) );
  XNOR2_X1 RoundFunction_T1_U346 ( .A(RoundFunction_STATE1[50]), .B(
        RoundFunction_T1_n590), .ZN(RoundFunction_TMP3_1[14]) );
  XNOR2_X1 RoundFunction_T1_U345 ( .A(RoundFunction_STATE1[4]), .B(
        RoundFunction_T1_n585), .ZN(RoundFunction_TMP3_1[4]) );
  XNOR2_X1 RoundFunction_T1_U344 ( .A(RoundFunction_STATE1[49]), .B(
        RoundFunction_T1_n600), .ZN(RoundFunction_TMP3_1[13]) );
  XNOR2_X1 RoundFunction_T1_U343 ( .A(RoundFunction_STATE1[48]), .B(
        RoundFunction_T1_n589), .ZN(RoundFunction_TMP3_1[12]) );
  XNOR2_X1 RoundFunction_T1_U342 ( .A(RoundFunction_STATE1[47]), .B(
        RoundFunction_T1_n588), .ZN(RoundFunction_TMP3_1[131]) );
  XNOR2_X1 RoundFunction_T1_U341 ( .A(RoundFunction_STATE1[46]), .B(
        RoundFunction_T1_n587), .ZN(RoundFunction_TMP3_1[130]) );
  XNOR2_X1 RoundFunction_T1_U340 ( .A(RoundFunction_STATE1[45]), .B(
        RoundFunction_T1_n586), .ZN(RoundFunction_TMP3_1[129]) );
  XNOR2_X1 RoundFunction_T1_U339 ( .A(RoundFunction_STATE1[44]), .B(
        RoundFunction_T1_n585), .ZN(RoundFunction_TMP3_1[128]) );
  XNOR2_X1 RoundFunction_T1_U338 ( .A(RoundFunction_STATE1[43]), .B(
        RoundFunction_T1_n584), .ZN(RoundFunction_TMP3_1[135]) );
  XNOR2_X1 RoundFunction_T1_U337 ( .A(RoundFunction_STATE1[42]), .B(
        RoundFunction_T1_n583), .ZN(RoundFunction_TMP3_1[134]) );
  XNOR2_X1 RoundFunction_T1_U336 ( .A(RoundFunction_STATE1[41]), .B(
        RoundFunction_T1_n582), .ZN(RoundFunction_TMP3_1[133]) );
  XNOR2_X1 RoundFunction_T1_U335 ( .A(RoundFunction_STATE1[40]), .B(
        RoundFunction_T1_n581), .ZN(RoundFunction_TMP3_1[132]) );
  XNOR2_X1 RoundFunction_T1_U334 ( .A(RoundFunction_STATE1[3]), .B(
        RoundFunction_T1_n584), .ZN(RoundFunction_TMP3_1[3]) );
  XNOR2_X1 RoundFunction_T1_U333 ( .A(RoundFunction_STATE1[39]), .B(
        RoundFunction_T1_n580), .ZN(RoundFunction_TMP3_1[122]) );
  XNOR2_X1 RoundFunction_T1_U332 ( .A(RoundFunction_STATE1[38]), .B(
        RoundFunction_T1_n579), .ZN(RoundFunction_TMP3_1[121]) );
  XNOR2_X1 RoundFunction_T1_U331 ( .A(RoundFunction_STATE1[37]), .B(
        RoundFunction_T1_n578), .ZN(RoundFunction_TMP3_1[120]) );
  XNOR2_X1 RoundFunction_T1_U330 ( .A(RoundFunction_STATE1[36]), .B(
        RoundFunction_T1_n577), .ZN(RoundFunction_TMP3_1[127]) );
  XNOR2_X1 RoundFunction_T1_U329 ( .A(RoundFunction_STATE1[35]), .B(
        RoundFunction_T1_n576), .ZN(RoundFunction_TMP3_1[126]) );
  XNOR2_X1 RoundFunction_T1_U328 ( .A(RoundFunction_STATE1[34]), .B(
        RoundFunction_T1_n575), .ZN(RoundFunction_TMP3_1[125]) );
  XNOR2_X1 RoundFunction_T1_U327 ( .A(RoundFunction_STATE1[33]), .B(
        RoundFunction_T1_n574), .ZN(RoundFunction_TMP3_1[124]) );
  XNOR2_X1 RoundFunction_T1_U326 ( .A(RoundFunction_STATE1[32]), .B(
        RoundFunction_T1_n573), .ZN(RoundFunction_TMP3_1[123]) );
  XNOR2_X1 RoundFunction_T1_U325 ( .A(RoundFunction_STATE1[31]), .B(
        RoundFunction_T1_n572), .ZN(RoundFunction_TMP3_1[43]) );
  XNOR2_X1 RoundFunction_T1_U324 ( .A(RoundFunction_STATE1[30]), .B(
        RoundFunction_T1_n571), .ZN(RoundFunction_TMP3_1[42]) );
  XNOR2_X1 RoundFunction_T1_U323 ( .A(RoundFunction_STATE1[2]), .B(
        RoundFunction_T1_n583), .ZN(RoundFunction_TMP3_1[2]) );
  XNOR2_X1 RoundFunction_T1_U322 ( .A(RoundFunction_STATE1[29]), .B(
        RoundFunction_T1_n570), .ZN(RoundFunction_TMP3_1[41]) );
  XNOR2_X1 RoundFunction_T1_U321 ( .A(RoundFunction_STATE1[28]), .B(
        RoundFunction_T1_n569), .ZN(RoundFunction_TMP3_1[40]) );
  XNOR2_X1 RoundFunction_T1_U320 ( .A(RoundFunction_STATE1[27]), .B(
        RoundFunction_T1_n568), .ZN(RoundFunction_TMP3_1[47]) );
  XNOR2_X1 RoundFunction_T1_U319 ( .A(RoundFunction_STATE1[26]), .B(
        RoundFunction_T1_n567), .ZN(RoundFunction_TMP3_1[46]) );
  XNOR2_X1 RoundFunction_T1_U318 ( .A(RoundFunction_STATE1[25]), .B(
        RoundFunction_T1_n566), .ZN(RoundFunction_TMP3_1[45]) );
  XNOR2_X1 RoundFunction_T1_U317 ( .A(RoundFunction_STATE1[24]), .B(
        RoundFunction_T1_n565), .ZN(RoundFunction_TMP3_1[44]) );
  XNOR2_X1 RoundFunction_T1_U316 ( .A(RoundFunction_STATE1[23]), .B(
        RoundFunction_T1_n564), .ZN(RoundFunction_TMP3_1[165]) );
  XNOR2_X1 RoundFunction_T1_U315 ( .A(RoundFunction_STATE1[22]), .B(
        RoundFunction_T1_n563), .ZN(RoundFunction_TMP3_1[164]) );
  XNOR2_X1 RoundFunction_T1_U314 ( .A(RoundFunction_STATE1[21]), .B(
        RoundFunction_T1_n562), .ZN(RoundFunction_TMP3_1[163]) );
  XNOR2_X1 RoundFunction_T1_U313 ( .A(RoundFunction_STATE1[20]), .B(
        RoundFunction_T1_n561), .ZN(RoundFunction_TMP3_1[162]) );
  XNOR2_X1 RoundFunction_T1_U312 ( .A(RoundFunction_STATE1[1]), .B(
        RoundFunction_T1_n582), .ZN(RoundFunction_TMP3_1[1]) );
  XNOR2_X1 RoundFunction_T1_U311 ( .A(RoundFunction_STATE1[19]), .B(
        RoundFunction_T1_n599), .ZN(RoundFunction_TMP3_1[161]) );
  XNOR2_X1 RoundFunction_T1_U310 ( .A(RoundFunction_STATE1[199]), .B(
        RoundFunction_T1_n580), .ZN(RoundFunction_TMP3_1[37]) );
  XNOR2_X1 RoundFunction_T1_U309 ( .A(RoundFunction_STATE1[198]), .B(
        RoundFunction_T1_n579), .ZN(RoundFunction_TMP3_1[36]) );
  XNOR2_X1 RoundFunction_T1_U308 ( .A(RoundFunction_STATE1[197]), .B(
        RoundFunction_T1_n578), .ZN(RoundFunction_TMP3_1[35]) );
  XNOR2_X1 RoundFunction_T1_U307 ( .A(RoundFunction_STATE1[196]), .B(
        RoundFunction_T1_n577), .ZN(RoundFunction_TMP3_1[34]) );
  XNOR2_X1 RoundFunction_T1_U306 ( .A(RoundFunction_STATE1[195]), .B(
        RoundFunction_T1_n576), .ZN(RoundFunction_TMP3_1[33]) );
  XNOR2_X1 RoundFunction_T1_U305 ( .A(RoundFunction_STATE1[194]), .B(
        RoundFunction_T1_n575), .ZN(RoundFunction_TMP3_1[32]) );
  XNOR2_X1 RoundFunction_T1_U304 ( .A(RoundFunction_STATE1[193]), .B(
        RoundFunction_T1_n574), .ZN(RoundFunction_TMP3_1[39]) );
  XNOR2_X1 RoundFunction_T1_U303 ( .A(RoundFunction_STATE1[192]), .B(
        RoundFunction_T1_n573), .ZN(RoundFunction_TMP3_1[38]) );
  XNOR2_X1 RoundFunction_T1_U302 ( .A(RoundFunction_STATE1[191]), .B(
        RoundFunction_T1_n572), .ZN(RoundFunction_TMP3_1[159]) );
  XNOR2_X1 RoundFunction_T1_U301 ( .A(RoundFunction_STATE1[190]), .B(
        RoundFunction_T1_n571), .ZN(RoundFunction_TMP3_1[158]) );
  XNOR2_X1 RoundFunction_T1_U300 ( .A(RoundFunction_STATE1[18]), .B(
        RoundFunction_T1_n598), .ZN(RoundFunction_TMP3_1[160]) );
  XNOR2_X1 RoundFunction_T1_U299 ( .A(RoundFunction_STATE1[189]), .B(
        RoundFunction_T1_n570), .ZN(RoundFunction_TMP3_1[157]) );
  XNOR2_X1 RoundFunction_T1_U298 ( .A(RoundFunction_STATE1[188]), .B(
        RoundFunction_T1_n569), .ZN(RoundFunction_TMP3_1[156]) );
  XNOR2_X1 RoundFunction_T1_U297 ( .A(RoundFunction_STATE1[187]), .B(
        RoundFunction_T1_n568), .ZN(RoundFunction_TMP3_1[155]) );
  XNOR2_X1 RoundFunction_T1_U296 ( .A(RoundFunction_STATE1[186]), .B(
        RoundFunction_T1_n567), .ZN(RoundFunction_TMP3_1[154]) );
  XNOR2_X1 RoundFunction_T1_U295 ( .A(RoundFunction_STATE1[185]), .B(
        RoundFunction_T1_n566), .ZN(RoundFunction_TMP3_1[153]) );
  XNOR2_X1 RoundFunction_T1_U294 ( .A(RoundFunction_STATE1[184]), .B(
        RoundFunction_T1_n565), .ZN(RoundFunction_TMP3_1[152]) );
  XNOR2_X1 RoundFunction_T1_U293 ( .A(RoundFunction_STATE1[183]), .B(
        RoundFunction_T1_n564), .ZN(RoundFunction_TMP3_1[76]) );
  XNOR2_X1 RoundFunction_T1_U292 ( .A(RoundFunction_STATE1[182]), .B(
        RoundFunction_T1_n563), .ZN(RoundFunction_TMP3_1[75]) );
  XNOR2_X1 RoundFunction_T1_U291 ( .A(RoundFunction_STATE1[181]), .B(
        RoundFunction_T1_n562), .ZN(RoundFunction_TMP3_1[74]) );
  XNOR2_X1 RoundFunction_T1_U290 ( .A(RoundFunction_STATE1[180]), .B(
        RoundFunction_T1_n561), .ZN(RoundFunction_TMP3_1[73]) );
  XNOR2_X1 RoundFunction_T1_U289 ( .A(RoundFunction_STATE1[17]), .B(
        RoundFunction_T1_n597), .ZN(RoundFunction_TMP3_1[167]) );
  XNOR2_X1 RoundFunction_T1_U288 ( .A(RoundFunction_STATE1[179]), .B(
        RoundFunction_T1_n599), .ZN(RoundFunction_TMP3_1[72]) );
  XNOR2_X1 RoundFunction_T1_U287 ( .A(RoundFunction_STATE1[178]), .B(
        RoundFunction_T1_n598), .ZN(RoundFunction_TMP3_1[79]) );
  XNOR2_X1 RoundFunction_T1_U286 ( .A(RoundFunction_STATE1[177]), .B(
        RoundFunction_T1_n597), .ZN(RoundFunction_TMP3_1[78]) );
  XNOR2_X1 RoundFunction_T1_U285 ( .A(RoundFunction_STATE1[176]), .B(
        RoundFunction_T1_n596), .ZN(RoundFunction_TMP3_1[77]) );
  XNOR2_X1 RoundFunction_T1_U284 ( .A(RoundFunction_STATE1[175]), .B(
        RoundFunction_T1_n595), .ZN(RoundFunction_TMP3_1[193]) );
  XNOR2_X1 RoundFunction_T1_U283 ( .A(RoundFunction_STATE1[174]), .B(
        RoundFunction_T1_n594), .ZN(RoundFunction_TMP3_1[192]) );
  XNOR2_X1 RoundFunction_T1_U282 ( .A(RoundFunction_STATE1[173]), .B(
        RoundFunction_T1_n593), .ZN(RoundFunction_TMP3_1[199]) );
  XNOR2_X1 RoundFunction_T1_U281 ( .A(RoundFunction_STATE1[172]), .B(
        RoundFunction_T1_n592), .ZN(RoundFunction_TMP3_1[198]) );
  XNOR2_X1 RoundFunction_T1_U280 ( .A(RoundFunction_STATE1[171]), .B(
        RoundFunction_T1_n591), .ZN(RoundFunction_TMP3_1[197]) );
  XNOR2_X1 RoundFunction_T1_U279 ( .A(RoundFunction_STATE1[170]), .B(
        RoundFunction_T1_n590), .ZN(RoundFunction_TMP3_1[196]) );
  XNOR2_X1 RoundFunction_T1_U278 ( .A(RoundFunction_STATE1[16]), .B(
        RoundFunction_T1_n596), .ZN(RoundFunction_TMP3_1[166]) );
  XNOR2_X1 RoundFunction_T1_U277 ( .A(RoundFunction_STATE1[169]), .B(
        RoundFunction_T1_n600), .ZN(RoundFunction_TMP3_1[195]) );
  XNOR2_X1 RoundFunction_T1_U276 ( .A(RoundFunction_STATE1[168]), .B(
        RoundFunction_T1_n589), .ZN(RoundFunction_TMP3_1[194]) );
  XNOR2_X1 RoundFunction_T1_U275 ( .A(RoundFunction_STATE1[167]), .B(
        RoundFunction_T1_n588), .ZN(RoundFunction_TMP3_1[113]) );
  XNOR2_X1 RoundFunction_T1_U274 ( .A(RoundFunction_STATE1[166]), .B(
        RoundFunction_T1_n587), .ZN(RoundFunction_TMP3_1[112]) );
  XNOR2_X1 RoundFunction_T1_U273 ( .A(RoundFunction_STATE1[165]), .B(
        RoundFunction_T1_n586), .ZN(RoundFunction_TMP3_1[119]) );
  XNOR2_X1 RoundFunction_T1_U272 ( .A(RoundFunction_STATE1[164]), .B(
        RoundFunction_T1_n585), .ZN(RoundFunction_TMP3_1[118]) );
  XNOR2_X1 RoundFunction_T1_U271 ( .A(RoundFunction_STATE1[163]), .B(
        RoundFunction_T1_n584), .ZN(RoundFunction_TMP3_1[117]) );
  XNOR2_X1 RoundFunction_T1_U270 ( .A(RoundFunction_STATE1[162]), .B(
        RoundFunction_T1_n583), .ZN(RoundFunction_TMP3_1[116]) );
  XNOR2_X1 RoundFunction_T1_U269 ( .A(RoundFunction_STATE1[161]), .B(
        RoundFunction_T1_n582), .ZN(RoundFunction_TMP3_1[115]) );
  XNOR2_X1 RoundFunction_T1_U268 ( .A(RoundFunction_STATE1[160]), .B(
        RoundFunction_T1_n581), .ZN(RoundFunction_TMP3_1[114]) );
  XNOR2_X1 RoundFunction_T1_U267 ( .A(RoundFunction_STATE1[15]), .B(
        RoundFunction_T1_n595), .ZN(RoundFunction_TMP3_1[80]) );
  XNOR2_X1 RoundFunction_T1_U266 ( .A(RoundFunction_STATE1[159]), .B(
        RoundFunction_T1_n580), .ZN(RoundFunction_TMP3_1[111]) );
  XNOR2_X1 RoundFunction_T1_U265 ( .A(RoundFunction_STATE1[158]), .B(
        RoundFunction_T1_n579), .ZN(RoundFunction_TMP3_1[110]) );
  XNOR2_X1 RoundFunction_T1_U264 ( .A(RoundFunction_STATE1[157]), .B(
        RoundFunction_T1_n578), .ZN(RoundFunction_TMP3_1[109]) );
  XNOR2_X1 RoundFunction_T1_U263 ( .A(RoundFunction_STATE1[156]), .B(
        RoundFunction_T1_n577), .ZN(RoundFunction_TMP3_1[108]) );
  XNOR2_X1 RoundFunction_T1_U262 ( .A(RoundFunction_STATE1[155]), .B(
        RoundFunction_T1_n576), .ZN(RoundFunction_TMP3_1[107]) );
  XNOR2_X1 RoundFunction_T1_U261 ( .A(RoundFunction_STATE1[154]), .B(
        RoundFunction_T1_n575), .ZN(RoundFunction_TMP3_1[106]) );
  XNOR2_X1 RoundFunction_T1_U260 ( .A(RoundFunction_STATE1[153]), .B(
        RoundFunction_T1_n574), .ZN(RoundFunction_TMP3_1[105]) );
  XNOR2_X1 RoundFunction_T1_U259 ( .A(RoundFunction_STATE1[152]), .B(
        RoundFunction_T1_n573), .ZN(RoundFunction_TMP3_1[104]) );
  XNOR2_X1 RoundFunction_T1_U258 ( .A(RoundFunction_STATE1[151]), .B(
        RoundFunction_T1_n572), .ZN(RoundFunction_TMP3_1[28]) );
  XNOR2_X1 RoundFunction_T1_U257 ( .A(RoundFunction_STATE1[150]), .B(
        RoundFunction_T1_n571), .ZN(RoundFunction_TMP3_1[27]) );
  XNOR2_X1 RoundFunction_T1_U256 ( .A(RoundFunction_STATE1[14]), .B(
        RoundFunction_T1_n594), .ZN(RoundFunction_TMP3_1[87]) );
  XNOR2_X1 RoundFunction_T1_U255 ( .A(RoundFunction_STATE1[149]), .B(
        RoundFunction_T1_n570), .ZN(RoundFunction_TMP3_1[26]) );
  XNOR2_X1 RoundFunction_T1_U254 ( .A(RoundFunction_STATE1[148]), .B(
        RoundFunction_T1_n569), .ZN(RoundFunction_TMP3_1[25]) );
  XNOR2_X1 RoundFunction_T1_U253 ( .A(RoundFunction_STATE1[147]), .B(
        RoundFunction_T1_n568), .ZN(RoundFunction_TMP3_1[24]) );
  XNOR2_X1 RoundFunction_T1_U252 ( .A(RoundFunction_STATE1[146]), .B(
        RoundFunction_T1_n567), .ZN(RoundFunction_TMP3_1[31]) );
  XNOR2_X1 RoundFunction_T1_U251 ( .A(RoundFunction_STATE1[145]), .B(
        RoundFunction_T1_n566), .ZN(RoundFunction_TMP3_1[30]) );
  XNOR2_X1 RoundFunction_T1_U250 ( .A(RoundFunction_STATE1[144]), .B(
        RoundFunction_T1_n565), .ZN(RoundFunction_TMP3_1[29]) );
  XNOR2_X1 RoundFunction_T1_U249 ( .A(RoundFunction_STATE1[143]), .B(
        RoundFunction_T1_n564), .ZN(RoundFunction_TMP3_1[150]) );
  XNOR2_X1 RoundFunction_T1_U248 ( .A(RoundFunction_STATE1[142]), .B(
        RoundFunction_T1_n563), .ZN(RoundFunction_TMP3_1[149]) );
  XNOR2_X1 RoundFunction_T1_U247 ( .A(RoundFunction_STATE1[141]), .B(
        RoundFunction_T1_n562), .ZN(RoundFunction_TMP3_1[148]) );
  XNOR2_X1 RoundFunction_T1_U246 ( .A(RoundFunction_STATE1[140]), .B(
        RoundFunction_T1_n561), .ZN(RoundFunction_TMP3_1[147]) );
  XNOR2_X1 RoundFunction_T1_U245 ( .A(RoundFunction_STATE1[13]), .B(
        RoundFunction_T1_n593), .ZN(RoundFunction_TMP3_1[86]) );
  XNOR2_X1 RoundFunction_T1_U244 ( .A(RoundFunction_STATE1[139]), .B(
        RoundFunction_T1_n599), .ZN(RoundFunction_TMP3_1[146]) );
  XNOR2_X1 RoundFunction_T1_U243 ( .A(RoundFunction_T1_n560), .B(
        RoundFunction_T1_n559), .ZN(RoundFunction_T1_n599) );
  XNOR2_X1 RoundFunction_T1_U242 ( .A(RoundFunction_STATE1[138]), .B(
        RoundFunction_T1_n598), .ZN(RoundFunction_TMP3_1[145]) );
  XNOR2_X1 RoundFunction_T1_U241 ( .A(RoundFunction_T1_n558), .B(
        RoundFunction_T1_n557), .ZN(RoundFunction_T1_n598) );
  XNOR2_X1 RoundFunction_T1_U240 ( .A(RoundFunction_STATE1[137]), .B(
        RoundFunction_T1_n597), .ZN(RoundFunction_TMP3_1[144]) );
  XNOR2_X1 RoundFunction_T1_U239 ( .A(RoundFunction_T1_n556), .B(
        RoundFunction_T1_n555), .ZN(RoundFunction_T1_n597) );
  XNOR2_X1 RoundFunction_T1_U238 ( .A(RoundFunction_STATE1[136]), .B(
        RoundFunction_T1_n596), .ZN(RoundFunction_TMP3_1[151]) );
  XNOR2_X1 RoundFunction_T1_U237 ( .A(RoundFunction_T1_n554), .B(
        RoundFunction_T1_n553), .ZN(RoundFunction_T1_n596) );
  XNOR2_X1 RoundFunction_T1_U236 ( .A(RoundFunction_STATE1[135]), .B(
        RoundFunction_T1_n595), .ZN(RoundFunction_TMP3_1[68]) );
  XNOR2_X1 RoundFunction_T1_U235 ( .A(RoundFunction_T1_n552), .B(
        RoundFunction_T1_n551), .ZN(RoundFunction_T1_n595) );
  XNOR2_X1 RoundFunction_T1_U234 ( .A(RoundFunction_STATE1[134]), .B(
        RoundFunction_T1_n594), .ZN(RoundFunction_TMP3_1[67]) );
  XNOR2_X1 RoundFunction_T1_U233 ( .A(RoundFunction_T1_n550), .B(
        RoundFunction_T1_n549), .ZN(RoundFunction_T1_n594) );
  XNOR2_X1 RoundFunction_T1_U232 ( .A(RoundFunction_STATE1[133]), .B(
        RoundFunction_T1_n593), .ZN(RoundFunction_TMP3_1[66]) );
  XNOR2_X1 RoundFunction_T1_U231 ( .A(RoundFunction_T1_n548), .B(
        RoundFunction_T1_n547), .ZN(RoundFunction_T1_n593) );
  XNOR2_X1 RoundFunction_T1_U230 ( .A(RoundFunction_STATE1[132]), .B(
        RoundFunction_T1_n592), .ZN(RoundFunction_TMP3_1[65]) );
  XNOR2_X1 RoundFunction_T1_U229 ( .A(RoundFunction_STATE1[131]), .B(
        RoundFunction_T1_n591), .ZN(RoundFunction_TMP3_1[64]) );
  XNOR2_X1 RoundFunction_T1_U228 ( .A(RoundFunction_STATE1[130]), .B(
        RoundFunction_T1_n590), .ZN(RoundFunction_TMP3_1[71]) );
  XNOR2_X1 RoundFunction_T1_U227 ( .A(RoundFunction_STATE1[12]), .B(
        RoundFunction_T1_n592), .ZN(RoundFunction_TMP3_1[85]) );
  XNOR2_X1 RoundFunction_T1_U226 ( .A(RoundFunction_T1_n546), .B(
        RoundFunction_T1_n545), .ZN(RoundFunction_T1_n592) );
  XNOR2_X1 RoundFunction_T1_U225 ( .A(RoundFunction_STATE1[129]), .B(
        RoundFunction_T1_n600), .ZN(RoundFunction_TMP3_1[70]) );
  XNOR2_X1 RoundFunction_T1_U224 ( .A(RoundFunction_T1_n544), .B(
        RoundFunction_T1_n543), .ZN(RoundFunction_T1_n600) );
  XNOR2_X1 RoundFunction_T1_U223 ( .A(RoundFunction_STATE1[128]), .B(
        RoundFunction_T1_n589), .ZN(RoundFunction_TMP3_1[69]) );
  XNOR2_X1 RoundFunction_T1_U222 ( .A(RoundFunction_T1_n542), .B(
        RoundFunction_T1_n541), .ZN(RoundFunction_T1_n589) );
  XNOR2_X1 RoundFunction_T1_U221 ( .A(RoundFunction_STATE1[127]), .B(
        RoundFunction_T1_n588), .ZN(RoundFunction_TMP3_1[184]) );
  XNOR2_X1 RoundFunction_T1_U220 ( .A(RoundFunction_T1_n540), .B(
        RoundFunction_T1_n539), .ZN(RoundFunction_T1_n588) );
  XNOR2_X1 RoundFunction_T1_U219 ( .A(RoundFunction_STATE1[126]), .B(
        RoundFunction_T1_n587), .ZN(RoundFunction_TMP3_1[191]) );
  XNOR2_X1 RoundFunction_T1_U218 ( .A(RoundFunction_T1_n538), .B(
        RoundFunction_T1_n537), .ZN(RoundFunction_T1_n587) );
  XNOR2_X1 RoundFunction_T1_U217 ( .A(RoundFunction_STATE1[125]), .B(
        RoundFunction_T1_n586), .ZN(RoundFunction_TMP3_1[190]) );
  XNOR2_X1 RoundFunction_T1_U216 ( .A(RoundFunction_T1_n536), .B(
        RoundFunction_T1_n535), .ZN(RoundFunction_T1_n586) );
  XNOR2_X1 RoundFunction_T1_U215 ( .A(RoundFunction_STATE1[124]), .B(
        RoundFunction_T1_n585), .ZN(RoundFunction_TMP3_1[189]) );
  XNOR2_X1 RoundFunction_T1_U214 ( .A(RoundFunction_T1_n534), .B(
        RoundFunction_T1_n559), .ZN(RoundFunction_T1_n585) );
  XOR2_X1 RoundFunction_T1_U213 ( .A(RoundFunction_STATE1[11]), .B(
        RoundFunction_T1_n533), .Z(RoundFunction_T1_n559) );
  XNOR2_X1 RoundFunction_T1_U212 ( .A(RoundFunction_T1_n532), .B(
        RoundFunction_T1_n531), .ZN(RoundFunction_T1_n533) );
  XNOR2_X1 RoundFunction_T1_U211 ( .A(RoundFunction_STATE1[51]), .B(
        RoundFunction_STATE1[91]), .ZN(RoundFunction_T1_n531) );
  XOR2_X1 RoundFunction_T1_U210 ( .A(RoundFunction_STATE1[131]), .B(
        RoundFunction_STATE1[171]), .Z(RoundFunction_T1_n532) );
  XNOR2_X1 RoundFunction_T1_U209 ( .A(RoundFunction_STATE1[123]), .B(
        RoundFunction_T1_n584), .ZN(RoundFunction_TMP3_1[188]) );
  XNOR2_X1 RoundFunction_T1_U208 ( .A(RoundFunction_T1_n530), .B(
        RoundFunction_T1_n557), .ZN(RoundFunction_T1_n584) );
  XOR2_X1 RoundFunction_T1_U207 ( .A(RoundFunction_STATE1[10]), .B(
        RoundFunction_T1_n529), .Z(RoundFunction_T1_n557) );
  XNOR2_X1 RoundFunction_T1_U206 ( .A(RoundFunction_T1_n528), .B(
        RoundFunction_T1_n527), .ZN(RoundFunction_T1_n529) );
  XNOR2_X1 RoundFunction_T1_U205 ( .A(RoundFunction_STATE1[50]), .B(
        RoundFunction_STATE1[90]), .ZN(RoundFunction_T1_n527) );
  XOR2_X1 RoundFunction_T1_U204 ( .A(RoundFunction_STATE1[130]), .B(
        RoundFunction_STATE1[170]), .Z(RoundFunction_T1_n528) );
  XNOR2_X1 RoundFunction_T1_U203 ( .A(RoundFunction_STATE1[122]), .B(
        RoundFunction_T1_n583), .ZN(RoundFunction_TMP3_1[187]) );
  XNOR2_X1 RoundFunction_T1_U202 ( .A(RoundFunction_T1_n526), .B(
        RoundFunction_T1_n555), .ZN(RoundFunction_T1_n583) );
  XOR2_X1 RoundFunction_T1_U201 ( .A(RoundFunction_STATE1[89]), .B(
        RoundFunction_T1_n525), .Z(RoundFunction_T1_n555) );
  XNOR2_X1 RoundFunction_T1_U200 ( .A(RoundFunction_T1_n524), .B(
        RoundFunction_T1_n523), .ZN(RoundFunction_T1_n525) );
  XNOR2_X1 RoundFunction_T1_U199 ( .A(RoundFunction_STATE1[129]), .B(
        RoundFunction_STATE1[49]), .ZN(RoundFunction_T1_n523) );
  XOR2_X1 RoundFunction_T1_U198 ( .A(RoundFunction_STATE1[169]), .B(
        RoundFunction_STATE1[9]), .Z(RoundFunction_T1_n524) );
  XNOR2_X1 RoundFunction_T1_U197 ( .A(RoundFunction_STATE1[121]), .B(
        RoundFunction_T1_n582), .ZN(RoundFunction_TMP3_1[186]) );
  XNOR2_X1 RoundFunction_T1_U196 ( .A(RoundFunction_T1_n522), .B(
        RoundFunction_T1_n553), .ZN(RoundFunction_T1_n582) );
  XOR2_X1 RoundFunction_T1_U195 ( .A(RoundFunction_STATE1[128]), .B(
        RoundFunction_T1_n521), .Z(RoundFunction_T1_n553) );
  XNOR2_X1 RoundFunction_T1_U194 ( .A(RoundFunction_T1_n520), .B(
        RoundFunction_T1_n519), .ZN(RoundFunction_T1_n521) );
  XNOR2_X1 RoundFunction_T1_U193 ( .A(RoundFunction_STATE1[48]), .B(
        RoundFunction_STATE1[8]), .ZN(RoundFunction_T1_n519) );
  XOR2_X1 RoundFunction_T1_U192 ( .A(RoundFunction_STATE1[88]), .B(
        RoundFunction_STATE1[168]), .Z(RoundFunction_T1_n520) );
  XNOR2_X1 RoundFunction_T1_U191 ( .A(RoundFunction_STATE1[120]), .B(
        RoundFunction_T1_n581), .ZN(RoundFunction_TMP3_1[185]) );
  XNOR2_X1 RoundFunction_T1_U190 ( .A(RoundFunction_STATE1[11]), .B(
        RoundFunction_T1_n591), .ZN(RoundFunction_TMP3_1[84]) );
  XNOR2_X1 RoundFunction_T1_U189 ( .A(RoundFunction_T1_n518), .B(
        RoundFunction_T1_n517), .ZN(RoundFunction_T1_n591) );
  XNOR2_X1 RoundFunction_T1_U188 ( .A(RoundFunction_STATE1[119]), .B(
        RoundFunction_T1_n580), .ZN(RoundFunction_TMP3_1[182]) );
  XNOR2_X1 RoundFunction_T1_U187 ( .A(RoundFunction_T1_n554), .B(
        RoundFunction_T1_n549), .ZN(RoundFunction_T1_n580) );
  XOR2_X1 RoundFunction_T1_U186 ( .A(RoundFunction_STATE1[126]), .B(
        RoundFunction_T1_n516), .Z(RoundFunction_T1_n549) );
  XNOR2_X1 RoundFunction_T1_U185 ( .A(RoundFunction_T1_n515), .B(
        RoundFunction_T1_n514), .ZN(RoundFunction_T1_n516) );
  XNOR2_X1 RoundFunction_T1_U184 ( .A(RoundFunction_STATE1[46]), .B(
        RoundFunction_STATE1[86]), .ZN(RoundFunction_T1_n514) );
  XOR2_X1 RoundFunction_T1_U183 ( .A(RoundFunction_STATE1[6]), .B(
        RoundFunction_STATE1[166]), .Z(RoundFunction_T1_n515) );
  XOR2_X1 RoundFunction_T1_U182 ( .A(RoundFunction_STATE1[111]), .B(
        RoundFunction_T1_n513), .Z(RoundFunction_T1_n554) );
  XNOR2_X1 RoundFunction_T1_U181 ( .A(RoundFunction_T1_n512), .B(
        RoundFunction_T1_n511), .ZN(RoundFunction_T1_n513) );
  XNOR2_X1 RoundFunction_T1_U180 ( .A(RoundFunction_STATE1[31]), .B(
        RoundFunction_STATE1[71]), .ZN(RoundFunction_T1_n511) );
  XOR2_X1 RoundFunction_T1_U179 ( .A(RoundFunction_STATE1[151]), .B(
        RoundFunction_STATE1[191]), .Z(RoundFunction_T1_n512) );
  XNOR2_X1 RoundFunction_T1_U178 ( .A(RoundFunction_STATE1[118]), .B(
        RoundFunction_T1_n579), .ZN(RoundFunction_TMP3_1[181]) );
  XNOR2_X1 RoundFunction_T1_U177 ( .A(RoundFunction_T1_n510), .B(
        RoundFunction_T1_n547), .ZN(RoundFunction_T1_n579) );
  XOR2_X1 RoundFunction_T1_U176 ( .A(RoundFunction_STATE1[125]), .B(
        RoundFunction_T1_n509), .Z(RoundFunction_T1_n547) );
  XNOR2_X1 RoundFunction_T1_U175 ( .A(RoundFunction_T1_n508), .B(
        RoundFunction_T1_n507), .ZN(RoundFunction_T1_n509) );
  XNOR2_X1 RoundFunction_T1_U174 ( .A(RoundFunction_STATE1[45]), .B(
        RoundFunction_STATE1[85]), .ZN(RoundFunction_T1_n507) );
  XOR2_X1 RoundFunction_T1_U173 ( .A(RoundFunction_STATE1[5]), .B(
        RoundFunction_STATE1[165]), .Z(RoundFunction_T1_n508) );
  XNOR2_X1 RoundFunction_T1_U172 ( .A(RoundFunction_STATE1[117]), .B(
        RoundFunction_T1_n578), .ZN(RoundFunction_TMP3_1[180]) );
  XNOR2_X1 RoundFunction_T1_U171 ( .A(RoundFunction_T1_n506), .B(
        RoundFunction_T1_n545), .ZN(RoundFunction_T1_n578) );
  XOR2_X1 RoundFunction_T1_U170 ( .A(RoundFunction_STATE1[124]), .B(
        RoundFunction_T1_n505), .Z(RoundFunction_T1_n545) );
  XNOR2_X1 RoundFunction_T1_U169 ( .A(RoundFunction_T1_n504), .B(
        RoundFunction_T1_n503), .ZN(RoundFunction_T1_n505) );
  XNOR2_X1 RoundFunction_T1_U168 ( .A(RoundFunction_STATE1[44]), .B(
        RoundFunction_STATE1[84]), .ZN(RoundFunction_T1_n503) );
  XOR2_X1 RoundFunction_T1_U167 ( .A(RoundFunction_STATE1[4]), .B(
        RoundFunction_STATE1[164]), .Z(RoundFunction_T1_n504) );
  XNOR2_X1 RoundFunction_T1_U166 ( .A(RoundFunction_STATE1[116]), .B(
        RoundFunction_T1_n577), .ZN(RoundFunction_TMP3_1[179]) );
  XNOR2_X1 RoundFunction_T1_U165 ( .A(RoundFunction_T1_n502), .B(
        RoundFunction_T1_n517), .ZN(RoundFunction_T1_n577) );
  XOR2_X1 RoundFunction_T1_U164 ( .A(RoundFunction_STATE1[123]), .B(
        RoundFunction_T1_n501), .Z(RoundFunction_T1_n517) );
  XNOR2_X1 RoundFunction_T1_U163 ( .A(RoundFunction_T1_n500), .B(
        RoundFunction_T1_n499), .ZN(RoundFunction_T1_n501) );
  XNOR2_X1 RoundFunction_T1_U162 ( .A(RoundFunction_STATE1[3]), .B(
        RoundFunction_STATE1[83]), .ZN(RoundFunction_T1_n499) );
  XOR2_X1 RoundFunction_T1_U161 ( .A(RoundFunction_STATE1[43]), .B(
        RoundFunction_STATE1[163]), .Z(RoundFunction_T1_n500) );
  XNOR2_X1 RoundFunction_T1_U160 ( .A(RoundFunction_STATE1[115]), .B(
        RoundFunction_T1_n576), .ZN(RoundFunction_TMP3_1[178]) );
  XNOR2_X1 RoundFunction_T1_U159 ( .A(RoundFunction_T1_n498), .B(
        RoundFunction_T1_n497), .ZN(RoundFunction_T1_n576) );
  XNOR2_X1 RoundFunction_T1_U158 ( .A(RoundFunction_STATE1[114]), .B(
        RoundFunction_T1_n575), .ZN(RoundFunction_TMP3_1[177]) );
  XNOR2_X1 RoundFunction_T1_U157 ( .A(RoundFunction_T1_n543), .B(
        RoundFunction_T1_n560), .ZN(RoundFunction_T1_n575) );
  XOR2_X1 RoundFunction_T1_U156 ( .A(RoundFunction_STATE1[106]), .B(
        RoundFunction_T1_n496), .Z(RoundFunction_T1_n560) );
  XNOR2_X1 RoundFunction_T1_U155 ( .A(RoundFunction_T1_n495), .B(
        RoundFunction_T1_n494), .ZN(RoundFunction_T1_n496) );
  XNOR2_X1 RoundFunction_T1_U154 ( .A(RoundFunction_STATE1[26]), .B(
        RoundFunction_STATE1[66]), .ZN(RoundFunction_T1_n494) );
  XOR2_X1 RoundFunction_T1_U153 ( .A(RoundFunction_STATE1[146]), .B(
        RoundFunction_STATE1[186]), .Z(RoundFunction_T1_n495) );
  XOR2_X1 RoundFunction_T1_U152 ( .A(RoundFunction_STATE1[121]), .B(
        RoundFunction_T1_n493), .Z(RoundFunction_T1_n543) );
  XNOR2_X1 RoundFunction_T1_U151 ( .A(RoundFunction_T1_n492), .B(
        RoundFunction_T1_n491), .ZN(RoundFunction_T1_n493) );
  XNOR2_X1 RoundFunction_T1_U150 ( .A(RoundFunction_STATE1[1]), .B(
        RoundFunction_STATE1[81]), .ZN(RoundFunction_T1_n491) );
  XOR2_X1 RoundFunction_T1_U149 ( .A(RoundFunction_STATE1[41]), .B(
        RoundFunction_STATE1[161]), .Z(RoundFunction_T1_n492) );
  XNOR2_X1 RoundFunction_T1_U148 ( .A(RoundFunction_STATE1[113]), .B(
        RoundFunction_T1_n574), .ZN(RoundFunction_TMP3_1[176]) );
  XNOR2_X1 RoundFunction_T1_U147 ( .A(RoundFunction_T1_n558), .B(
        RoundFunction_T1_n541), .ZN(RoundFunction_T1_n574) );
  XOR2_X1 RoundFunction_T1_U146 ( .A(RoundFunction_STATE1[0]), .B(
        RoundFunction_T1_n490), .Z(RoundFunction_T1_n541) );
  XNOR2_X1 RoundFunction_T1_U145 ( .A(RoundFunction_T1_n489), .B(
        RoundFunction_T1_n488), .ZN(RoundFunction_T1_n490) );
  XNOR2_X1 RoundFunction_T1_U144 ( .A(RoundFunction_STATE1[40]), .B(
        RoundFunction_STATE1[80]), .ZN(RoundFunction_T1_n488) );
  XOR2_X1 RoundFunction_T1_U143 ( .A(RoundFunction_STATE1[120]), .B(
        RoundFunction_STATE1[160]), .Z(RoundFunction_T1_n489) );
  XOR2_X1 RoundFunction_T1_U142 ( .A(RoundFunction_STATE1[105]), .B(
        RoundFunction_T1_n487), .Z(RoundFunction_T1_n558) );
  XNOR2_X1 RoundFunction_T1_U141 ( .A(RoundFunction_T1_n486), .B(
        RoundFunction_T1_n485), .ZN(RoundFunction_T1_n487) );
  XNOR2_X1 RoundFunction_T1_U140 ( .A(RoundFunction_STATE1[25]), .B(
        RoundFunction_STATE1[65]), .ZN(RoundFunction_T1_n485) );
  XOR2_X1 RoundFunction_T1_U139 ( .A(RoundFunction_STATE1[145]), .B(
        RoundFunction_STATE1[185]), .Z(RoundFunction_T1_n486) );
  XNOR2_X1 RoundFunction_T1_U138 ( .A(RoundFunction_STATE1[112]), .B(
        RoundFunction_T1_n573), .ZN(RoundFunction_TMP3_1[183]) );
  XNOR2_X1 RoundFunction_T1_U137 ( .A(RoundFunction_T1_n556), .B(
        RoundFunction_T1_n551), .ZN(RoundFunction_T1_n573) );
  XOR2_X1 RoundFunction_T1_U136 ( .A(RoundFunction_STATE1[127]), .B(
        RoundFunction_T1_n484), .Z(RoundFunction_T1_n551) );
  XNOR2_X1 RoundFunction_T1_U135 ( .A(RoundFunction_T1_n483), .B(
        RoundFunction_T1_n482), .ZN(RoundFunction_T1_n484) );
  XNOR2_X1 RoundFunction_T1_U134 ( .A(RoundFunction_STATE1[47]), .B(
        RoundFunction_STATE1[87]), .ZN(RoundFunction_T1_n482) );
  XOR2_X1 RoundFunction_T1_U133 ( .A(RoundFunction_STATE1[7]), .B(
        RoundFunction_STATE1[167]), .Z(RoundFunction_T1_n483) );
  XOR2_X1 RoundFunction_T1_U132 ( .A(RoundFunction_STATE1[104]), .B(
        RoundFunction_T1_n481), .Z(RoundFunction_T1_n556) );
  XNOR2_X1 RoundFunction_T1_U131 ( .A(RoundFunction_T1_n480), .B(
        RoundFunction_T1_n479), .ZN(RoundFunction_T1_n481) );
  XNOR2_X1 RoundFunction_T1_U130 ( .A(RoundFunction_STATE1[24]), .B(
        RoundFunction_STATE1[64]), .ZN(RoundFunction_T1_n479) );
  XOR2_X1 RoundFunction_T1_U129 ( .A(RoundFunction_STATE1[144]), .B(
        RoundFunction_STATE1[184]), .Z(RoundFunction_T1_n480) );
  XNOR2_X1 RoundFunction_T1_U128 ( .A(RoundFunction_STATE1[111]), .B(
        RoundFunction_T1_n572), .ZN(RoundFunction_TMP3_1[96]) );
  XNOR2_X1 RoundFunction_T1_U127 ( .A(RoundFunction_T1_n542), .B(
        RoundFunction_T1_n537), .ZN(RoundFunction_T1_n572) );
  XOR2_X1 RoundFunction_T1_U126 ( .A(RoundFunction_STATE1[118]), .B(
        RoundFunction_T1_n478), .Z(RoundFunction_T1_n537) );
  XNOR2_X1 RoundFunction_T1_U125 ( .A(RoundFunction_T1_n477), .B(
        RoundFunction_T1_n476), .ZN(RoundFunction_T1_n478) );
  XNOR2_X1 RoundFunction_T1_U124 ( .A(RoundFunction_STATE1[198]), .B(
        RoundFunction_STATE1[78]), .ZN(RoundFunction_T1_n476) );
  XOR2_X1 RoundFunction_T1_U123 ( .A(RoundFunction_STATE1[38]), .B(
        RoundFunction_STATE1[158]), .Z(RoundFunction_T1_n477) );
  XOR2_X1 RoundFunction_T1_U122 ( .A(RoundFunction_STATE1[103]), .B(
        RoundFunction_T1_n475), .Z(RoundFunction_T1_n542) );
  XNOR2_X1 RoundFunction_T1_U121 ( .A(RoundFunction_T1_n474), .B(
        RoundFunction_T1_n473), .ZN(RoundFunction_T1_n475) );
  XNOR2_X1 RoundFunction_T1_U120 ( .A(RoundFunction_STATE1[23]), .B(
        RoundFunction_STATE1[63]), .ZN(RoundFunction_T1_n473) );
  XOR2_X1 RoundFunction_T1_U119 ( .A(RoundFunction_STATE1[143]), .B(
        RoundFunction_STATE1[183]), .Z(RoundFunction_T1_n474) );
  XNOR2_X1 RoundFunction_T1_U118 ( .A(RoundFunction_STATE1[110]), .B(
        RoundFunction_T1_n571), .ZN(RoundFunction_TMP3_1[103]) );
  XNOR2_X1 RoundFunction_T1_U117 ( .A(RoundFunction_T1_n552), .B(
        RoundFunction_T1_n535), .ZN(RoundFunction_T1_n571) );
  XOR2_X1 RoundFunction_T1_U116 ( .A(RoundFunction_STATE1[117]), .B(
        RoundFunction_T1_n472), .Z(RoundFunction_T1_n535) );
  XNOR2_X1 RoundFunction_T1_U115 ( .A(RoundFunction_T1_n471), .B(
        RoundFunction_T1_n470), .ZN(RoundFunction_T1_n472) );
  XNOR2_X1 RoundFunction_T1_U114 ( .A(RoundFunction_STATE1[197]), .B(
        RoundFunction_STATE1[77]), .ZN(RoundFunction_T1_n470) );
  XOR2_X1 RoundFunction_T1_U113 ( .A(RoundFunction_STATE1[37]), .B(
        RoundFunction_STATE1[157]), .Z(RoundFunction_T1_n471) );
  XOR2_X1 RoundFunction_T1_U112 ( .A(RoundFunction_STATE1[102]), .B(
        RoundFunction_T1_n469), .Z(RoundFunction_T1_n552) );
  XNOR2_X1 RoundFunction_T1_U111 ( .A(RoundFunction_T1_n468), .B(
        RoundFunction_T1_n467), .ZN(RoundFunction_T1_n469) );
  XNOR2_X1 RoundFunction_T1_U110 ( .A(RoundFunction_STATE1[22]), .B(
        RoundFunction_STATE1[62]), .ZN(RoundFunction_T1_n467) );
  XOR2_X1 RoundFunction_T1_U109 ( .A(RoundFunction_STATE1[142]), .B(
        RoundFunction_STATE1[182]), .Z(RoundFunction_T1_n468) );
  XNOR2_X1 RoundFunction_T1_U108 ( .A(RoundFunction_STATE1[10]), .B(
        RoundFunction_T1_n590), .ZN(RoundFunction_TMP3_1[83]) );
  XNOR2_X1 RoundFunction_T1_U107 ( .A(RoundFunction_T1_n466), .B(
        RoundFunction_T1_n497), .ZN(RoundFunction_T1_n590) );
  XOR2_X1 RoundFunction_T1_U106 ( .A(RoundFunction_STATE1[122]), .B(
        RoundFunction_T1_n465), .Z(RoundFunction_T1_n497) );
  XNOR2_X1 RoundFunction_T1_U105 ( .A(RoundFunction_T1_n464), .B(
        RoundFunction_T1_n463), .ZN(RoundFunction_T1_n465) );
  XNOR2_X1 RoundFunction_T1_U104 ( .A(RoundFunction_STATE1[2]), .B(
        RoundFunction_STATE1[82]), .ZN(RoundFunction_T1_n463) );
  XOR2_X1 RoundFunction_T1_U103 ( .A(RoundFunction_STATE1[42]), .B(
        RoundFunction_STATE1[162]), .Z(RoundFunction_T1_n464) );
  XNOR2_X1 RoundFunction_T1_U102 ( .A(RoundFunction_STATE1[109]), .B(
        RoundFunction_T1_n570), .ZN(RoundFunction_TMP3_1[102]) );
  XNOR2_X1 RoundFunction_T1_U101 ( .A(RoundFunction_T1_n550), .B(
        RoundFunction_T1_n534), .ZN(RoundFunction_T1_n570) );
  XOR2_X1 RoundFunction_T1_U100 ( .A(RoundFunction_STATE1[116]), .B(
        RoundFunction_T1_n462), .Z(RoundFunction_T1_n534) );
  XNOR2_X1 RoundFunction_T1_U99 ( .A(RoundFunction_T1_n461), .B(
        RoundFunction_T1_n460), .ZN(RoundFunction_T1_n462) );
  XNOR2_X1 RoundFunction_T1_U98 ( .A(RoundFunction_STATE1[196]), .B(
        RoundFunction_STATE1[76]), .ZN(RoundFunction_T1_n460) );
  XOR2_X1 RoundFunction_T1_U97 ( .A(RoundFunction_STATE1[36]), .B(
        RoundFunction_STATE1[156]), .Z(RoundFunction_T1_n461) );
  XOR2_X1 RoundFunction_T1_U96 ( .A(RoundFunction_STATE1[101]), .B(
        RoundFunction_T1_n459), .Z(RoundFunction_T1_n550) );
  XNOR2_X1 RoundFunction_T1_U95 ( .A(RoundFunction_T1_n458), .B(
        RoundFunction_T1_n457), .ZN(RoundFunction_T1_n459) );
  XNOR2_X1 RoundFunction_T1_U94 ( .A(RoundFunction_STATE1[21]), .B(
        RoundFunction_STATE1[61]), .ZN(RoundFunction_T1_n457) );
  XOR2_X1 RoundFunction_T1_U93 ( .A(RoundFunction_STATE1[141]), .B(
        RoundFunction_STATE1[181]), .Z(RoundFunction_T1_n458) );
  XNOR2_X1 RoundFunction_T1_U92 ( .A(RoundFunction_STATE1[108]), .B(
        RoundFunction_T1_n569), .ZN(RoundFunction_TMP3_1[101]) );
  XNOR2_X1 RoundFunction_T1_U91 ( .A(RoundFunction_T1_n548), .B(
        RoundFunction_T1_n530), .ZN(RoundFunction_T1_n569) );
  XOR2_X1 RoundFunction_T1_U90 ( .A(RoundFunction_STATE1[115]), .B(
        RoundFunction_T1_n456), .Z(RoundFunction_T1_n530) );
  XNOR2_X1 RoundFunction_T1_U89 ( .A(RoundFunction_T1_n455), .B(
        RoundFunction_T1_n454), .ZN(RoundFunction_T1_n456) );
  XNOR2_X1 RoundFunction_T1_U88 ( .A(RoundFunction_STATE1[195]), .B(
        RoundFunction_STATE1[75]), .ZN(RoundFunction_T1_n454) );
  XOR2_X1 RoundFunction_T1_U87 ( .A(RoundFunction_STATE1[35]), .B(
        RoundFunction_STATE1[155]), .Z(RoundFunction_T1_n455) );
  XOR2_X1 RoundFunction_T1_U86 ( .A(RoundFunction_STATE1[100]), .B(
        RoundFunction_T1_n453), .Z(RoundFunction_T1_n548) );
  XNOR2_X1 RoundFunction_T1_U85 ( .A(RoundFunction_T1_n452), .B(
        RoundFunction_T1_n451), .ZN(RoundFunction_T1_n453) );
  XNOR2_X1 RoundFunction_T1_U84 ( .A(RoundFunction_STATE1[20]), .B(
        RoundFunction_STATE1[60]), .ZN(RoundFunction_T1_n451) );
  XOR2_X1 RoundFunction_T1_U83 ( .A(RoundFunction_STATE1[140]), .B(
        RoundFunction_STATE1[180]), .Z(RoundFunction_T1_n452) );
  XNOR2_X1 RoundFunction_T1_U82 ( .A(RoundFunction_STATE1[107]), .B(
        RoundFunction_T1_n568), .ZN(RoundFunction_TMP3_1[100]) );
  XNOR2_X1 RoundFunction_T1_U81 ( .A(RoundFunction_T1_n546), .B(
        RoundFunction_T1_n526), .ZN(RoundFunction_T1_n568) );
  XOR2_X1 RoundFunction_T1_U80 ( .A(RoundFunction_STATE1[114]), .B(
        RoundFunction_T1_n450), .Z(RoundFunction_T1_n526) );
  XNOR2_X1 RoundFunction_T1_U79 ( .A(RoundFunction_T1_n449), .B(
        RoundFunction_T1_n448), .ZN(RoundFunction_T1_n450) );
  XNOR2_X1 RoundFunction_T1_U78 ( .A(RoundFunction_STATE1[194]), .B(
        RoundFunction_STATE1[74]), .ZN(RoundFunction_T1_n448) );
  XOR2_X1 RoundFunction_T1_U77 ( .A(RoundFunction_STATE1[34]), .B(
        RoundFunction_STATE1[154]), .Z(RoundFunction_T1_n449) );
  XOR2_X1 RoundFunction_T1_U76 ( .A(RoundFunction_STATE1[59]), .B(
        RoundFunction_T1_n447), .Z(RoundFunction_T1_n546) );
  XNOR2_X1 RoundFunction_T1_U75 ( .A(RoundFunction_T1_n446), .B(
        RoundFunction_T1_n445), .ZN(RoundFunction_T1_n447) );
  XNOR2_X1 RoundFunction_T1_U74 ( .A(RoundFunction_STATE1[139]), .B(
        RoundFunction_STATE1[19]), .ZN(RoundFunction_T1_n445) );
  XOR2_X1 RoundFunction_T1_U73 ( .A(RoundFunction_STATE1[179]), .B(
        RoundFunction_STATE1[99]), .Z(RoundFunction_T1_n446) );
  XNOR2_X1 RoundFunction_T1_U72 ( .A(RoundFunction_STATE1[106]), .B(
        RoundFunction_T1_n567), .ZN(RoundFunction_TMP3_1[99]) );
  XNOR2_X1 RoundFunction_T1_U71 ( .A(RoundFunction_T1_n518), .B(
        RoundFunction_T1_n522), .ZN(RoundFunction_T1_n567) );
  XOR2_X1 RoundFunction_T1_U70 ( .A(RoundFunction_STATE1[113]), .B(
        RoundFunction_T1_n444), .Z(RoundFunction_T1_n522) );
  XNOR2_X1 RoundFunction_T1_U69 ( .A(RoundFunction_T1_n443), .B(
        RoundFunction_T1_n442), .ZN(RoundFunction_T1_n444) );
  XNOR2_X1 RoundFunction_T1_U68 ( .A(RoundFunction_STATE1[193]), .B(
        RoundFunction_STATE1[73]), .ZN(RoundFunction_T1_n442) );
  XOR2_X1 RoundFunction_T1_U67 ( .A(RoundFunction_STATE1[33]), .B(
        RoundFunction_STATE1[153]), .Z(RoundFunction_T1_n443) );
  XOR2_X1 RoundFunction_T1_U66 ( .A(RoundFunction_STATE1[58]), .B(
        RoundFunction_T1_n441), .Z(RoundFunction_T1_n518) );
  XNOR2_X1 RoundFunction_T1_U65 ( .A(RoundFunction_T1_n440), .B(
        RoundFunction_T1_n439), .ZN(RoundFunction_T1_n441) );
  XNOR2_X1 RoundFunction_T1_U64 ( .A(RoundFunction_STATE1[138]), .B(
        RoundFunction_STATE1[18]), .ZN(RoundFunction_T1_n439) );
  XOR2_X1 RoundFunction_T1_U63 ( .A(RoundFunction_STATE1[178]), .B(
        RoundFunction_STATE1[98]), .Z(RoundFunction_T1_n440) );
  XNOR2_X1 RoundFunction_T1_U62 ( .A(RoundFunction_STATE1[105]), .B(
        RoundFunction_T1_n566), .ZN(RoundFunction_TMP3_1[98]) );
  XNOR2_X1 RoundFunction_T1_U61 ( .A(RoundFunction_T1_n438), .B(
        RoundFunction_T1_n466), .ZN(RoundFunction_T1_n566) );
  XOR2_X1 RoundFunction_T1_U60 ( .A(RoundFunction_STATE1[57]), .B(
        RoundFunction_T1_n437), .Z(RoundFunction_T1_n466) );
  XNOR2_X1 RoundFunction_T1_U59 ( .A(RoundFunction_T1_n436), .B(
        RoundFunction_T1_n435), .ZN(RoundFunction_T1_n437) );
  XNOR2_X1 RoundFunction_T1_U58 ( .A(RoundFunction_STATE1[137]), .B(
        RoundFunction_STATE1[17]), .ZN(RoundFunction_T1_n435) );
  XOR2_X1 RoundFunction_T1_U57 ( .A(RoundFunction_STATE1[177]), .B(
        RoundFunction_STATE1[97]), .Z(RoundFunction_T1_n436) );
  XNOR2_X1 RoundFunction_T1_U56 ( .A(RoundFunction_STATE1[104]), .B(
        RoundFunction_T1_n565), .ZN(RoundFunction_TMP3_1[97]) );
  XNOR2_X1 RoundFunction_T1_U55 ( .A(RoundFunction_T1_n544), .B(
        RoundFunction_T1_n539), .ZN(RoundFunction_T1_n565) );
  XOR2_X1 RoundFunction_T1_U54 ( .A(RoundFunction_STATE1[119]), .B(
        RoundFunction_T1_n434), .Z(RoundFunction_T1_n539) );
  XNOR2_X1 RoundFunction_T1_U53 ( .A(RoundFunction_T1_n433), .B(
        RoundFunction_T1_n432), .ZN(RoundFunction_T1_n434) );
  XNOR2_X1 RoundFunction_T1_U52 ( .A(RoundFunction_STATE1[199]), .B(
        RoundFunction_STATE1[79]), .ZN(RoundFunction_T1_n432) );
  XOR2_X1 RoundFunction_T1_U51 ( .A(RoundFunction_STATE1[39]), .B(
        RoundFunction_STATE1[159]), .Z(RoundFunction_T1_n433) );
  XOR2_X1 RoundFunction_T1_U50 ( .A(RoundFunction_STATE1[136]), .B(
        RoundFunction_T1_n431), .Z(RoundFunction_T1_n544) );
  XNOR2_X1 RoundFunction_T1_U49 ( .A(RoundFunction_T1_n430), .B(
        RoundFunction_T1_n429), .ZN(RoundFunction_T1_n431) );
  XNOR2_X1 RoundFunction_T1_U48 ( .A(RoundFunction_STATE1[176]), .B(
        RoundFunction_STATE1[96]), .ZN(RoundFunction_T1_n429) );
  XOR2_X1 RoundFunction_T1_U47 ( .A(RoundFunction_STATE1[56]), .B(
        RoundFunction_STATE1[16]), .Z(RoundFunction_T1_n430) );
  XNOR2_X1 RoundFunction_T1_U46 ( .A(RoundFunction_STATE1[103]), .B(
        RoundFunction_T1_n564), .ZN(RoundFunction_TMP3_1[18]) );
  XNOR2_X1 RoundFunction_T1_U45 ( .A(RoundFunction_T1_n428), .B(
        RoundFunction_T1_n510), .ZN(RoundFunction_T1_n564) );
  XOR2_X1 RoundFunction_T1_U44 ( .A(RoundFunction_STATE1[110]), .B(
        RoundFunction_T1_n427), .Z(RoundFunction_T1_n510) );
  XNOR2_X1 RoundFunction_T1_U43 ( .A(RoundFunction_T1_n426), .B(
        RoundFunction_T1_n425), .ZN(RoundFunction_T1_n427) );
  XNOR2_X1 RoundFunction_T1_U42 ( .A(RoundFunction_STATE1[190]), .B(
        RoundFunction_STATE1[70]), .ZN(RoundFunction_T1_n425) );
  XOR2_X1 RoundFunction_T1_U41 ( .A(RoundFunction_STATE1[30]), .B(
        RoundFunction_STATE1[150]), .Z(RoundFunction_T1_n426) );
  XNOR2_X1 RoundFunction_T1_U40 ( .A(RoundFunction_STATE1[102]), .B(
        RoundFunction_T1_n563), .ZN(RoundFunction_TMP3_1[17]) );
  XNOR2_X1 RoundFunction_T1_U39 ( .A(RoundFunction_T1_n540), .B(
        RoundFunction_T1_n506), .ZN(RoundFunction_T1_n563) );
  XOR2_X1 RoundFunction_T1_U38 ( .A(RoundFunction_STATE1[109]), .B(
        RoundFunction_T1_n424), .Z(RoundFunction_T1_n506) );
  XNOR2_X1 RoundFunction_T1_U37 ( .A(RoundFunction_T1_n423), .B(
        RoundFunction_T1_n422), .ZN(RoundFunction_T1_n424) );
  XNOR2_X1 RoundFunction_T1_U36 ( .A(RoundFunction_STATE1[189]), .B(
        RoundFunction_STATE1[69]), .ZN(RoundFunction_T1_n422) );
  XOR2_X1 RoundFunction_T1_U35 ( .A(RoundFunction_STATE1[29]), .B(
        RoundFunction_STATE1[149]), .Z(RoundFunction_T1_n423) );
  XOR2_X1 RoundFunction_T1_U34 ( .A(RoundFunction_STATE1[54]), .B(
        RoundFunction_T1_n421), .Z(RoundFunction_T1_n540) );
  XNOR2_X1 RoundFunction_T1_U33 ( .A(RoundFunction_T1_n420), .B(
        RoundFunction_T1_n419), .ZN(RoundFunction_T1_n421) );
  XNOR2_X1 RoundFunction_T1_U32 ( .A(RoundFunction_STATE1[134]), .B(
        RoundFunction_STATE1[174]), .ZN(RoundFunction_T1_n419) );
  XOR2_X1 RoundFunction_T1_U31 ( .A(RoundFunction_STATE1[14]), .B(
        RoundFunction_STATE1[94]), .Z(RoundFunction_T1_n420) );
  XNOR2_X1 RoundFunction_T1_U30 ( .A(RoundFunction_STATE1[101]), .B(
        RoundFunction_T1_n562), .ZN(RoundFunction_TMP3_1[16]) );
  XNOR2_X1 RoundFunction_T1_U29 ( .A(RoundFunction_T1_n538), .B(
        RoundFunction_T1_n502), .ZN(RoundFunction_T1_n562) );
  XOR2_X1 RoundFunction_T1_U28 ( .A(RoundFunction_STATE1[108]), .B(
        RoundFunction_T1_n418), .Z(RoundFunction_T1_n502) );
  XNOR2_X1 RoundFunction_T1_U27 ( .A(RoundFunction_T1_n417), .B(
        RoundFunction_T1_n416), .ZN(RoundFunction_T1_n418) );
  XNOR2_X1 RoundFunction_T1_U26 ( .A(RoundFunction_STATE1[188]), .B(
        RoundFunction_STATE1[68]), .ZN(RoundFunction_T1_n416) );
  XOR2_X1 RoundFunction_T1_U25 ( .A(RoundFunction_STATE1[28]), .B(
        RoundFunction_STATE1[148]), .Z(RoundFunction_T1_n417) );
  XOR2_X1 RoundFunction_T1_U24 ( .A(RoundFunction_STATE1[53]), .B(
        RoundFunction_T1_n415), .Z(RoundFunction_T1_n538) );
  XNOR2_X1 RoundFunction_T1_U23 ( .A(RoundFunction_T1_n414), .B(
        RoundFunction_T1_n413), .ZN(RoundFunction_T1_n415) );
  XNOR2_X1 RoundFunction_T1_U22 ( .A(RoundFunction_STATE1[133]), .B(
        RoundFunction_STATE1[173]), .ZN(RoundFunction_T1_n413) );
  XOR2_X1 RoundFunction_T1_U21 ( .A(RoundFunction_STATE1[13]), .B(
        RoundFunction_STATE1[93]), .Z(RoundFunction_T1_n414) );
  XNOR2_X1 RoundFunction_T1_U20 ( .A(RoundFunction_STATE1[100]), .B(
        RoundFunction_T1_n561), .ZN(RoundFunction_TMP3_1[23]) );
  XNOR2_X1 RoundFunction_T1_U19 ( .A(RoundFunction_T1_n536), .B(
        RoundFunction_T1_n498), .ZN(RoundFunction_T1_n561) );
  XOR2_X1 RoundFunction_T1_U18 ( .A(RoundFunction_STATE1[107]), .B(
        RoundFunction_T1_n412), .Z(RoundFunction_T1_n498) );
  XNOR2_X1 RoundFunction_T1_U17 ( .A(RoundFunction_T1_n411), .B(
        RoundFunction_T1_n410), .ZN(RoundFunction_T1_n412) );
  XNOR2_X1 RoundFunction_T1_U16 ( .A(RoundFunction_STATE1[187]), .B(
        RoundFunction_STATE1[67]), .ZN(RoundFunction_T1_n410) );
  XOR2_X1 RoundFunction_T1_U15 ( .A(RoundFunction_STATE1[27]), .B(
        RoundFunction_STATE1[147]), .Z(RoundFunction_T1_n411) );
  XOR2_X1 RoundFunction_T1_U14 ( .A(RoundFunction_STATE1[52]), .B(
        RoundFunction_T1_n409), .Z(RoundFunction_T1_n536) );
  XNOR2_X1 RoundFunction_T1_U13 ( .A(RoundFunction_T1_n408), .B(
        RoundFunction_T1_n407), .ZN(RoundFunction_T1_n409) );
  XNOR2_X1 RoundFunction_T1_U12 ( .A(RoundFunction_STATE1[12]), .B(
        RoundFunction_STATE1[172]), .ZN(RoundFunction_T1_n407) );
  XOR2_X1 RoundFunction_T1_U11 ( .A(RoundFunction_STATE1[132]), .B(
        RoundFunction_STATE1[92]), .Z(RoundFunction_T1_n408) );
  XNOR2_X1 RoundFunction_T1_U10 ( .A(RoundFunction_STATE1[0]), .B(
        RoundFunction_T1_n581), .ZN(RoundFunction_TMP3_1[0]) );
  XNOR2_X1 RoundFunction_T1_U9 ( .A(RoundFunction_T1_n438), .B(
        RoundFunction_T1_n428), .ZN(RoundFunction_T1_n581) );
  XOR2_X1 RoundFunction_T1_U8 ( .A(RoundFunction_STATE1[55]), .B(
        RoundFunction_T1_n406), .Z(RoundFunction_T1_n428) );
  XNOR2_X1 RoundFunction_T1_U7 ( .A(RoundFunction_T1_n405), .B(
        RoundFunction_T1_n404), .ZN(RoundFunction_T1_n406) );
  XNOR2_X1 RoundFunction_T1_U6 ( .A(RoundFunction_STATE1[135]), .B(
        RoundFunction_STATE1[175]), .ZN(RoundFunction_T1_n404) );
  XOR2_X1 RoundFunction_T1_U5 ( .A(RoundFunction_STATE1[15]), .B(
        RoundFunction_STATE1[95]), .Z(RoundFunction_T1_n405) );
  XOR2_X1 RoundFunction_T1_U4 ( .A(RoundFunction_STATE1[112]), .B(
        RoundFunction_T1_n403), .Z(RoundFunction_T1_n438) );
  XNOR2_X1 RoundFunction_T1_U3 ( .A(RoundFunction_T1_n402), .B(
        RoundFunction_T1_n401), .ZN(RoundFunction_T1_n403) );
  XNOR2_X1 RoundFunction_T1_U2 ( .A(RoundFunction_STATE1[192]), .B(
        RoundFunction_STATE1[72]), .ZN(RoundFunction_T1_n401) );
  XOR2_X1 RoundFunction_T1_U1 ( .A(RoundFunction_STATE1[32]), .B(
        RoundFunction_STATE1[152]), .Z(RoundFunction_T1_n402) );
  XOR2_X1 RoundFunction_I1_U8 ( .A(CONST[7]), .B(RoundFunction_TMP4_1[7]), .Z(
        RESULT1[199]) );
  XOR2_X1 RoundFunction_I1_U7 ( .A(1'b0), .B(RoundFunction_TMP4_1[6]), .Z(
        RESULT1[198]) );
  XOR2_X1 RoundFunction_I1_U6 ( .A(1'b0), .B(RoundFunction_TMP4_1[5]), .Z(
        RESULT1[197]) );
  XOR2_X1 RoundFunction_I1_U5 ( .A(1'b0), .B(RoundFunction_TMP4_1[4]), .Z(
        RESULT1[196]) );
  XOR2_X1 RoundFunction_I1_U4 ( .A(CONST[3]), .B(RoundFunction_TMP4_1[3]), .Z(
        RESULT1[195]) );
  XOR2_X1 RoundFunction_I1_U3 ( .A(1'b0), .B(RoundFunction_TMP4_1[2]), .Z(
        RESULT1[194]) );
  XOR2_X1 RoundFunction_I1_U2 ( .A(CONST[1]), .B(RoundFunction_TMP4_1[1]), .Z(
        RESULT1[193]) );
  XOR2_X1 RoundFunction_I1_U1 ( .A(CONST[0]), .B(RoundFunction_TMP4_1[0]), .Z(
        RESULT1[192]) );
  XNOR2_X1 RoundFunction_T2_U400 ( .A(RoundFunction_STATE2[9]), .B(
        RoundFunction_T2_n600), .ZN(RoundFunction_TMP3_2[82]) );
  XNOR2_X1 RoundFunction_T2_U399 ( .A(RoundFunction_STATE2[99]), .B(
        RoundFunction_T2_n599), .ZN(RoundFunction_TMP3_2[22]) );
  XNOR2_X1 RoundFunction_T2_U398 ( .A(RoundFunction_STATE2[98]), .B(
        RoundFunction_T2_n598), .ZN(RoundFunction_TMP3_2[21]) );
  XNOR2_X1 RoundFunction_T2_U397 ( .A(RoundFunction_STATE2[97]), .B(
        RoundFunction_T2_n597), .ZN(RoundFunction_TMP3_2[20]) );
  XNOR2_X1 RoundFunction_T2_U396 ( .A(RoundFunction_STATE2[96]), .B(
        RoundFunction_T2_n596), .ZN(RoundFunction_TMP3_2[19]) );
  XNOR2_X1 RoundFunction_T2_U395 ( .A(RoundFunction_STATE2[95]), .B(
        RoundFunction_T2_n595), .ZN(RoundFunction_TMP3_2[137]) );
  XNOR2_X1 RoundFunction_T2_U394 ( .A(RoundFunction_STATE2[94]), .B(
        RoundFunction_T2_n594), .ZN(RoundFunction_TMP3_2[136]) );
  XNOR2_X1 RoundFunction_T2_U393 ( .A(RoundFunction_STATE2[93]), .B(
        RoundFunction_T2_n593), .ZN(RoundFunction_TMP3_2[143]) );
  XNOR2_X1 RoundFunction_T2_U392 ( .A(RoundFunction_STATE2[92]), .B(
        RoundFunction_T2_n592), .ZN(RoundFunction_TMP3_2[142]) );
  XNOR2_X1 RoundFunction_T2_U391 ( .A(RoundFunction_STATE2[91]), .B(
        RoundFunction_T2_n591), .ZN(RoundFunction_TMP3_2[141]) );
  XNOR2_X1 RoundFunction_T2_U390 ( .A(RoundFunction_STATE2[90]), .B(
        RoundFunction_T2_n590), .ZN(RoundFunction_TMP3_2[140]) );
  XNOR2_X1 RoundFunction_T2_U389 ( .A(RoundFunction_STATE2[8]), .B(
        RoundFunction_T2_n589), .ZN(RoundFunction_TMP3_2[81]) );
  XNOR2_X1 RoundFunction_T2_U388 ( .A(RoundFunction_STATE2[89]), .B(
        RoundFunction_T2_n600), .ZN(RoundFunction_TMP3_2[139]) );
  XNOR2_X1 RoundFunction_T2_U387 ( .A(RoundFunction_STATE2[88]), .B(
        RoundFunction_T2_n589), .ZN(RoundFunction_TMP3_2[138]) );
  XNOR2_X1 RoundFunction_T2_U386 ( .A(RoundFunction_STATE2[87]), .B(
        RoundFunction_T2_n588), .ZN(RoundFunction_TMP3_2[58]) );
  XNOR2_X1 RoundFunction_T2_U385 ( .A(RoundFunction_STATE2[86]), .B(
        RoundFunction_T2_n587), .ZN(RoundFunction_TMP3_2[57]) );
  XNOR2_X1 RoundFunction_T2_U384 ( .A(RoundFunction_STATE2[85]), .B(
        RoundFunction_T2_n586), .ZN(RoundFunction_TMP3_2[56]) );
  XNOR2_X1 RoundFunction_T2_U383 ( .A(RoundFunction_STATE2[84]), .B(
        RoundFunction_T2_n585), .ZN(RoundFunction_TMP3_2[63]) );
  XNOR2_X1 RoundFunction_T2_U382 ( .A(RoundFunction_STATE2[83]), .B(
        RoundFunction_T2_n584), .ZN(RoundFunction_TMP3_2[62]) );
  XNOR2_X1 RoundFunction_T2_U381 ( .A(RoundFunction_STATE2[82]), .B(
        RoundFunction_T2_n583), .ZN(RoundFunction_TMP3_2[61]) );
  XNOR2_X1 RoundFunction_T2_U380 ( .A(RoundFunction_STATE2[81]), .B(
        RoundFunction_T2_n582), .ZN(RoundFunction_TMP3_2[60]) );
  XNOR2_X1 RoundFunction_T2_U379 ( .A(RoundFunction_STATE2[80]), .B(
        RoundFunction_T2_n581), .ZN(RoundFunction_TMP3_2[59]) );
  XNOR2_X1 RoundFunction_T2_U378 ( .A(RoundFunction_STATE2[7]), .B(
        RoundFunction_T2_n588), .ZN(RoundFunction_TMP3_2[7]) );
  XNOR2_X1 RoundFunction_T2_U377 ( .A(RoundFunction_STATE2[79]), .B(
        RoundFunction_T2_n580), .ZN(RoundFunction_TMP3_2[51]) );
  XNOR2_X1 RoundFunction_T2_U376 ( .A(RoundFunction_STATE2[78]), .B(
        RoundFunction_T2_n579), .ZN(RoundFunction_TMP3_2[50]) );
  XNOR2_X1 RoundFunction_T2_U375 ( .A(RoundFunction_STATE2[77]), .B(
        RoundFunction_T2_n578), .ZN(RoundFunction_TMP3_2[49]) );
  XNOR2_X1 RoundFunction_T2_U374 ( .A(RoundFunction_STATE2[76]), .B(
        RoundFunction_T2_n577), .ZN(RoundFunction_TMP3_2[48]) );
  XNOR2_X1 RoundFunction_T2_U373 ( .A(RoundFunction_STATE2[75]), .B(
        RoundFunction_T2_n576), .ZN(RoundFunction_TMP3_2[55]) );
  XNOR2_X1 RoundFunction_T2_U372 ( .A(RoundFunction_STATE2[74]), .B(
        RoundFunction_T2_n575), .ZN(RoundFunction_TMP3_2[54]) );
  XNOR2_X1 RoundFunction_T2_U371 ( .A(RoundFunction_STATE2[73]), .B(
        RoundFunction_T2_n574), .ZN(RoundFunction_TMP3_2[53]) );
  XNOR2_X1 RoundFunction_T2_U370 ( .A(RoundFunction_STATE2[72]), .B(
        RoundFunction_T2_n573), .ZN(RoundFunction_TMP3_2[52]) );
  XNOR2_X1 RoundFunction_T2_U369 ( .A(RoundFunction_STATE2[71]), .B(
        RoundFunction_T2_n572), .ZN(RoundFunction_TMP3_2[174]) );
  XNOR2_X1 RoundFunction_T2_U368 ( .A(RoundFunction_STATE2[70]), .B(
        RoundFunction_T2_n571), .ZN(RoundFunction_TMP3_2[173]) );
  XNOR2_X1 RoundFunction_T2_U367 ( .A(RoundFunction_STATE2[6]), .B(
        RoundFunction_T2_n587), .ZN(RoundFunction_TMP3_2[6]) );
  XNOR2_X1 RoundFunction_T2_U366 ( .A(RoundFunction_STATE2[69]), .B(
        RoundFunction_T2_n570), .ZN(RoundFunction_TMP3_2[172]) );
  XNOR2_X1 RoundFunction_T2_U365 ( .A(RoundFunction_STATE2[68]), .B(
        RoundFunction_T2_n569), .ZN(RoundFunction_TMP3_2[171]) );
  XNOR2_X1 RoundFunction_T2_U364 ( .A(RoundFunction_STATE2[67]), .B(
        RoundFunction_T2_n568), .ZN(RoundFunction_TMP3_2[170]) );
  XNOR2_X1 RoundFunction_T2_U363 ( .A(RoundFunction_STATE2[66]), .B(
        RoundFunction_T2_n567), .ZN(RoundFunction_TMP3_2[169]) );
  XNOR2_X1 RoundFunction_T2_U362 ( .A(RoundFunction_STATE2[65]), .B(
        RoundFunction_T2_n566), .ZN(RoundFunction_TMP3_2[168]) );
  XNOR2_X1 RoundFunction_T2_U361 ( .A(RoundFunction_STATE2[64]), .B(
        RoundFunction_T2_n565), .ZN(RoundFunction_TMP3_2[175]) );
  XNOR2_X1 RoundFunction_T2_U360 ( .A(RoundFunction_STATE2[63]), .B(
        RoundFunction_T2_n564), .ZN(RoundFunction_TMP3_2[93]) );
  XNOR2_X1 RoundFunction_T2_U359 ( .A(RoundFunction_STATE2[62]), .B(
        RoundFunction_T2_n563), .ZN(RoundFunction_TMP3_2[92]) );
  XNOR2_X1 RoundFunction_T2_U358 ( .A(RoundFunction_STATE2[61]), .B(
        RoundFunction_T2_n562), .ZN(RoundFunction_TMP3_2[91]) );
  XNOR2_X1 RoundFunction_T2_U357 ( .A(RoundFunction_STATE2[60]), .B(
        RoundFunction_T2_n561), .ZN(RoundFunction_TMP3_2[90]) );
  XNOR2_X1 RoundFunction_T2_U356 ( .A(RoundFunction_STATE2[5]), .B(
        RoundFunction_T2_n586), .ZN(RoundFunction_TMP3_2[5]) );
  XNOR2_X1 RoundFunction_T2_U355 ( .A(RoundFunction_STATE2[59]), .B(
        RoundFunction_T2_n599), .ZN(RoundFunction_TMP3_2[89]) );
  XNOR2_X1 RoundFunction_T2_U354 ( .A(RoundFunction_STATE2[58]), .B(
        RoundFunction_T2_n598), .ZN(RoundFunction_TMP3_2[88]) );
  XNOR2_X1 RoundFunction_T2_U353 ( .A(RoundFunction_STATE2[57]), .B(
        RoundFunction_T2_n597), .ZN(RoundFunction_TMP3_2[95]) );
  XNOR2_X1 RoundFunction_T2_U352 ( .A(RoundFunction_STATE2[56]), .B(
        RoundFunction_T2_n596), .ZN(RoundFunction_TMP3_2[94]) );
  XNOR2_X1 RoundFunction_T2_U351 ( .A(RoundFunction_STATE2[55]), .B(
        RoundFunction_T2_n595), .ZN(RoundFunction_TMP3_2[11]) );
  XNOR2_X1 RoundFunction_T2_U350 ( .A(RoundFunction_STATE2[54]), .B(
        RoundFunction_T2_n594), .ZN(RoundFunction_TMP3_2[10]) );
  XNOR2_X1 RoundFunction_T2_U349 ( .A(RoundFunction_STATE2[53]), .B(
        RoundFunction_T2_n593), .ZN(RoundFunction_TMP3_2[9]) );
  XNOR2_X1 RoundFunction_T2_U348 ( .A(RoundFunction_STATE2[52]), .B(
        RoundFunction_T2_n592), .ZN(RoundFunction_TMP3_2[8]) );
  XNOR2_X1 RoundFunction_T2_U347 ( .A(RoundFunction_STATE2[51]), .B(
        RoundFunction_T2_n591), .ZN(RoundFunction_TMP3_2[15]) );
  XNOR2_X1 RoundFunction_T2_U346 ( .A(RoundFunction_STATE2[50]), .B(
        RoundFunction_T2_n590), .ZN(RoundFunction_TMP3_2[14]) );
  XNOR2_X1 RoundFunction_T2_U345 ( .A(RoundFunction_STATE2[4]), .B(
        RoundFunction_T2_n585), .ZN(RoundFunction_TMP3_2[4]) );
  XNOR2_X1 RoundFunction_T2_U344 ( .A(RoundFunction_STATE2[49]), .B(
        RoundFunction_T2_n600), .ZN(RoundFunction_TMP3_2[13]) );
  XNOR2_X1 RoundFunction_T2_U343 ( .A(RoundFunction_STATE2[48]), .B(
        RoundFunction_T2_n589), .ZN(RoundFunction_TMP3_2[12]) );
  XNOR2_X1 RoundFunction_T2_U342 ( .A(RoundFunction_STATE2[47]), .B(
        RoundFunction_T2_n588), .ZN(RoundFunction_TMP3_2[131]) );
  XNOR2_X1 RoundFunction_T2_U341 ( .A(RoundFunction_STATE2[46]), .B(
        RoundFunction_T2_n587), .ZN(RoundFunction_TMP3_2[130]) );
  XNOR2_X1 RoundFunction_T2_U340 ( .A(RoundFunction_STATE2[45]), .B(
        RoundFunction_T2_n586), .ZN(RoundFunction_TMP3_2[129]) );
  XNOR2_X1 RoundFunction_T2_U339 ( .A(RoundFunction_STATE2[44]), .B(
        RoundFunction_T2_n585), .ZN(RoundFunction_TMP3_2[128]) );
  XNOR2_X1 RoundFunction_T2_U338 ( .A(RoundFunction_STATE2[43]), .B(
        RoundFunction_T2_n584), .ZN(RoundFunction_TMP3_2[135]) );
  XNOR2_X1 RoundFunction_T2_U337 ( .A(RoundFunction_STATE2[42]), .B(
        RoundFunction_T2_n583), .ZN(RoundFunction_TMP3_2[134]) );
  XNOR2_X1 RoundFunction_T2_U336 ( .A(RoundFunction_STATE2[41]), .B(
        RoundFunction_T2_n582), .ZN(RoundFunction_TMP3_2[133]) );
  XNOR2_X1 RoundFunction_T2_U335 ( .A(RoundFunction_STATE2[40]), .B(
        RoundFunction_T2_n581), .ZN(RoundFunction_TMP3_2[132]) );
  XNOR2_X1 RoundFunction_T2_U334 ( .A(RoundFunction_STATE2[3]), .B(
        RoundFunction_T2_n584), .ZN(RoundFunction_TMP3_2[3]) );
  XNOR2_X1 RoundFunction_T2_U333 ( .A(RoundFunction_STATE2[39]), .B(
        RoundFunction_T2_n580), .ZN(RoundFunction_TMP3_2[122]) );
  XNOR2_X1 RoundFunction_T2_U332 ( .A(RoundFunction_STATE2[38]), .B(
        RoundFunction_T2_n579), .ZN(RoundFunction_TMP3_2[121]) );
  XNOR2_X1 RoundFunction_T2_U331 ( .A(RoundFunction_STATE2[37]), .B(
        RoundFunction_T2_n578), .ZN(RoundFunction_TMP3_2[120]) );
  XNOR2_X1 RoundFunction_T2_U330 ( .A(RoundFunction_STATE2[36]), .B(
        RoundFunction_T2_n577), .ZN(RoundFunction_TMP3_2[127]) );
  XNOR2_X1 RoundFunction_T2_U329 ( .A(RoundFunction_STATE2[35]), .B(
        RoundFunction_T2_n576), .ZN(RoundFunction_TMP3_2[126]) );
  XNOR2_X1 RoundFunction_T2_U328 ( .A(RoundFunction_STATE2[34]), .B(
        RoundFunction_T2_n575), .ZN(RoundFunction_TMP3_2[125]) );
  XNOR2_X1 RoundFunction_T2_U327 ( .A(RoundFunction_STATE2[33]), .B(
        RoundFunction_T2_n574), .ZN(RoundFunction_TMP3_2[124]) );
  XNOR2_X1 RoundFunction_T2_U326 ( .A(RoundFunction_STATE2[32]), .B(
        RoundFunction_T2_n573), .ZN(RoundFunction_TMP3_2[123]) );
  XNOR2_X1 RoundFunction_T2_U325 ( .A(RoundFunction_STATE2[31]), .B(
        RoundFunction_T2_n572), .ZN(RoundFunction_TMP3_2[43]) );
  XNOR2_X1 RoundFunction_T2_U324 ( .A(RoundFunction_STATE2[30]), .B(
        RoundFunction_T2_n571), .ZN(RoundFunction_TMP3_2[42]) );
  XNOR2_X1 RoundFunction_T2_U323 ( .A(RoundFunction_STATE2[2]), .B(
        RoundFunction_T2_n583), .ZN(RoundFunction_TMP3_2[2]) );
  XNOR2_X1 RoundFunction_T2_U322 ( .A(RoundFunction_STATE2[29]), .B(
        RoundFunction_T2_n570), .ZN(RoundFunction_TMP3_2[41]) );
  XNOR2_X1 RoundFunction_T2_U321 ( .A(RoundFunction_STATE2[28]), .B(
        RoundFunction_T2_n569), .ZN(RoundFunction_TMP3_2[40]) );
  XNOR2_X1 RoundFunction_T2_U320 ( .A(RoundFunction_STATE2[27]), .B(
        RoundFunction_T2_n568), .ZN(RoundFunction_TMP3_2[47]) );
  XNOR2_X1 RoundFunction_T2_U319 ( .A(RoundFunction_STATE2[26]), .B(
        RoundFunction_T2_n567), .ZN(RoundFunction_TMP3_2[46]) );
  XNOR2_X1 RoundFunction_T2_U318 ( .A(RoundFunction_STATE2[25]), .B(
        RoundFunction_T2_n566), .ZN(RoundFunction_TMP3_2[45]) );
  XNOR2_X1 RoundFunction_T2_U317 ( .A(RoundFunction_STATE2[24]), .B(
        RoundFunction_T2_n565), .ZN(RoundFunction_TMP3_2[44]) );
  XNOR2_X1 RoundFunction_T2_U316 ( .A(RoundFunction_STATE2[23]), .B(
        RoundFunction_T2_n564), .ZN(RoundFunction_TMP3_2[165]) );
  XNOR2_X1 RoundFunction_T2_U315 ( .A(RoundFunction_STATE2[22]), .B(
        RoundFunction_T2_n563), .ZN(RoundFunction_TMP3_2[164]) );
  XNOR2_X1 RoundFunction_T2_U314 ( .A(RoundFunction_STATE2[21]), .B(
        RoundFunction_T2_n562), .ZN(RoundFunction_TMP3_2[163]) );
  XNOR2_X1 RoundFunction_T2_U313 ( .A(RoundFunction_STATE2[20]), .B(
        RoundFunction_T2_n561), .ZN(RoundFunction_TMP3_2[162]) );
  XNOR2_X1 RoundFunction_T2_U312 ( .A(RoundFunction_STATE2[1]), .B(
        RoundFunction_T2_n582), .ZN(RoundFunction_TMP3_2[1]) );
  XNOR2_X1 RoundFunction_T2_U311 ( .A(RoundFunction_STATE2[19]), .B(
        RoundFunction_T2_n599), .ZN(RoundFunction_TMP3_2[161]) );
  XNOR2_X1 RoundFunction_T2_U310 ( .A(RoundFunction_STATE2[199]), .B(
        RoundFunction_T2_n580), .ZN(RoundFunction_TMP3_2[37]) );
  XNOR2_X1 RoundFunction_T2_U309 ( .A(RoundFunction_STATE2[198]), .B(
        RoundFunction_T2_n579), .ZN(RoundFunction_TMP3_2[36]) );
  XNOR2_X1 RoundFunction_T2_U308 ( .A(RoundFunction_STATE2[197]), .B(
        RoundFunction_T2_n578), .ZN(RoundFunction_TMP3_2[35]) );
  XNOR2_X1 RoundFunction_T2_U307 ( .A(RoundFunction_STATE2[196]), .B(
        RoundFunction_T2_n577), .ZN(RoundFunction_TMP3_2[34]) );
  XNOR2_X1 RoundFunction_T2_U306 ( .A(RoundFunction_STATE2[195]), .B(
        RoundFunction_T2_n576), .ZN(RoundFunction_TMP3_2[33]) );
  XNOR2_X1 RoundFunction_T2_U305 ( .A(RoundFunction_STATE2[194]), .B(
        RoundFunction_T2_n575), .ZN(RoundFunction_TMP3_2[32]) );
  XNOR2_X1 RoundFunction_T2_U304 ( .A(RoundFunction_STATE2[193]), .B(
        RoundFunction_T2_n574), .ZN(RoundFunction_TMP3_2[39]) );
  XNOR2_X1 RoundFunction_T2_U303 ( .A(RoundFunction_STATE2[192]), .B(
        RoundFunction_T2_n573), .ZN(RoundFunction_TMP3_2[38]) );
  XNOR2_X1 RoundFunction_T2_U302 ( .A(RoundFunction_STATE2[191]), .B(
        RoundFunction_T2_n572), .ZN(RoundFunction_TMP3_2[159]) );
  XNOR2_X1 RoundFunction_T2_U301 ( .A(RoundFunction_STATE2[190]), .B(
        RoundFunction_T2_n571), .ZN(RoundFunction_TMP3_2[158]) );
  XNOR2_X1 RoundFunction_T2_U300 ( .A(RoundFunction_STATE2[18]), .B(
        RoundFunction_T2_n598), .ZN(RoundFunction_TMP3_2[160]) );
  XNOR2_X1 RoundFunction_T2_U299 ( .A(RoundFunction_STATE2[189]), .B(
        RoundFunction_T2_n570), .ZN(RoundFunction_TMP3_2[157]) );
  XNOR2_X1 RoundFunction_T2_U298 ( .A(RoundFunction_STATE2[188]), .B(
        RoundFunction_T2_n569), .ZN(RoundFunction_TMP3_2[156]) );
  XNOR2_X1 RoundFunction_T2_U297 ( .A(RoundFunction_STATE2[187]), .B(
        RoundFunction_T2_n568), .ZN(RoundFunction_TMP3_2[155]) );
  XNOR2_X1 RoundFunction_T2_U296 ( .A(RoundFunction_STATE2[186]), .B(
        RoundFunction_T2_n567), .ZN(RoundFunction_TMP3_2[154]) );
  XNOR2_X1 RoundFunction_T2_U295 ( .A(RoundFunction_STATE2[185]), .B(
        RoundFunction_T2_n566), .ZN(RoundFunction_TMP3_2[153]) );
  XNOR2_X1 RoundFunction_T2_U294 ( .A(RoundFunction_STATE2[184]), .B(
        RoundFunction_T2_n565), .ZN(RoundFunction_TMP3_2[152]) );
  XNOR2_X1 RoundFunction_T2_U293 ( .A(RoundFunction_STATE2[183]), .B(
        RoundFunction_T2_n564), .ZN(RoundFunction_TMP3_2[76]) );
  XNOR2_X1 RoundFunction_T2_U292 ( .A(RoundFunction_STATE2[182]), .B(
        RoundFunction_T2_n563), .ZN(RoundFunction_TMP3_2[75]) );
  XNOR2_X1 RoundFunction_T2_U291 ( .A(RoundFunction_STATE2[181]), .B(
        RoundFunction_T2_n562), .ZN(RoundFunction_TMP3_2[74]) );
  XNOR2_X1 RoundFunction_T2_U290 ( .A(RoundFunction_STATE2[180]), .B(
        RoundFunction_T2_n561), .ZN(RoundFunction_TMP3_2[73]) );
  XNOR2_X1 RoundFunction_T2_U289 ( .A(RoundFunction_STATE2[17]), .B(
        RoundFunction_T2_n597), .ZN(RoundFunction_TMP3_2[167]) );
  XNOR2_X1 RoundFunction_T2_U288 ( .A(RoundFunction_STATE2[179]), .B(
        RoundFunction_T2_n599), .ZN(RoundFunction_TMP3_2[72]) );
  XNOR2_X1 RoundFunction_T2_U287 ( .A(RoundFunction_STATE2[178]), .B(
        RoundFunction_T2_n598), .ZN(RoundFunction_TMP3_2[79]) );
  XNOR2_X1 RoundFunction_T2_U286 ( .A(RoundFunction_STATE2[177]), .B(
        RoundFunction_T2_n597), .ZN(RoundFunction_TMP3_2[78]) );
  XNOR2_X1 RoundFunction_T2_U285 ( .A(RoundFunction_STATE2[176]), .B(
        RoundFunction_T2_n596), .ZN(RoundFunction_TMP3_2[77]) );
  XNOR2_X1 RoundFunction_T2_U284 ( .A(RoundFunction_STATE2[175]), .B(
        RoundFunction_T2_n595), .ZN(RoundFunction_TMP3_2[193]) );
  XNOR2_X1 RoundFunction_T2_U283 ( .A(RoundFunction_STATE2[174]), .B(
        RoundFunction_T2_n594), .ZN(RoundFunction_TMP3_2[192]) );
  XNOR2_X1 RoundFunction_T2_U282 ( .A(RoundFunction_STATE2[173]), .B(
        RoundFunction_T2_n593), .ZN(RoundFunction_TMP3_2[199]) );
  XNOR2_X1 RoundFunction_T2_U281 ( .A(RoundFunction_STATE2[172]), .B(
        RoundFunction_T2_n592), .ZN(RoundFunction_TMP3_2[198]) );
  XNOR2_X1 RoundFunction_T2_U280 ( .A(RoundFunction_STATE2[171]), .B(
        RoundFunction_T2_n591), .ZN(RoundFunction_TMP3_2[197]) );
  XNOR2_X1 RoundFunction_T2_U279 ( .A(RoundFunction_STATE2[170]), .B(
        RoundFunction_T2_n590), .ZN(RoundFunction_TMP3_2[196]) );
  XNOR2_X1 RoundFunction_T2_U278 ( .A(RoundFunction_STATE2[16]), .B(
        RoundFunction_T2_n596), .ZN(RoundFunction_TMP3_2[166]) );
  XNOR2_X1 RoundFunction_T2_U277 ( .A(RoundFunction_STATE2[169]), .B(
        RoundFunction_T2_n600), .ZN(RoundFunction_TMP3_2[195]) );
  XNOR2_X1 RoundFunction_T2_U276 ( .A(RoundFunction_STATE2[168]), .B(
        RoundFunction_T2_n589), .ZN(RoundFunction_TMP3_2[194]) );
  XNOR2_X1 RoundFunction_T2_U275 ( .A(RoundFunction_STATE2[167]), .B(
        RoundFunction_T2_n588), .ZN(RoundFunction_TMP3_2[113]) );
  XNOR2_X1 RoundFunction_T2_U274 ( .A(RoundFunction_STATE2[166]), .B(
        RoundFunction_T2_n587), .ZN(RoundFunction_TMP3_2[112]) );
  XNOR2_X1 RoundFunction_T2_U273 ( .A(RoundFunction_STATE2[165]), .B(
        RoundFunction_T2_n586), .ZN(RoundFunction_TMP3_2[119]) );
  XNOR2_X1 RoundFunction_T2_U272 ( .A(RoundFunction_STATE2[164]), .B(
        RoundFunction_T2_n585), .ZN(RoundFunction_TMP3_2[118]) );
  XNOR2_X1 RoundFunction_T2_U271 ( .A(RoundFunction_STATE2[163]), .B(
        RoundFunction_T2_n584), .ZN(RoundFunction_TMP3_2[117]) );
  XNOR2_X1 RoundFunction_T2_U270 ( .A(RoundFunction_STATE2[162]), .B(
        RoundFunction_T2_n583), .ZN(RoundFunction_TMP3_2[116]) );
  XNOR2_X1 RoundFunction_T2_U269 ( .A(RoundFunction_STATE2[161]), .B(
        RoundFunction_T2_n582), .ZN(RoundFunction_TMP3_2[115]) );
  XNOR2_X1 RoundFunction_T2_U268 ( .A(RoundFunction_STATE2[160]), .B(
        RoundFunction_T2_n581), .ZN(RoundFunction_TMP3_2[114]) );
  XNOR2_X1 RoundFunction_T2_U267 ( .A(RoundFunction_STATE2[15]), .B(
        RoundFunction_T2_n595), .ZN(RoundFunction_TMP3_2[80]) );
  XNOR2_X1 RoundFunction_T2_U266 ( .A(RoundFunction_STATE2[159]), .B(
        RoundFunction_T2_n580), .ZN(RoundFunction_TMP3_2[111]) );
  XNOR2_X1 RoundFunction_T2_U265 ( .A(RoundFunction_STATE2[158]), .B(
        RoundFunction_T2_n579), .ZN(RoundFunction_TMP3_2[110]) );
  XNOR2_X1 RoundFunction_T2_U264 ( .A(RoundFunction_STATE2[157]), .B(
        RoundFunction_T2_n578), .ZN(RoundFunction_TMP3_2[109]) );
  XNOR2_X1 RoundFunction_T2_U263 ( .A(RoundFunction_STATE2[156]), .B(
        RoundFunction_T2_n577), .ZN(RoundFunction_TMP3_2[108]) );
  XNOR2_X1 RoundFunction_T2_U262 ( .A(RoundFunction_STATE2[155]), .B(
        RoundFunction_T2_n576), .ZN(RoundFunction_TMP3_2[107]) );
  XNOR2_X1 RoundFunction_T2_U261 ( .A(RoundFunction_STATE2[154]), .B(
        RoundFunction_T2_n575), .ZN(RoundFunction_TMP3_2[106]) );
  XNOR2_X1 RoundFunction_T2_U260 ( .A(RoundFunction_STATE2[153]), .B(
        RoundFunction_T2_n574), .ZN(RoundFunction_TMP3_2[105]) );
  XNOR2_X1 RoundFunction_T2_U259 ( .A(RoundFunction_STATE2[152]), .B(
        RoundFunction_T2_n573), .ZN(RoundFunction_TMP3_2[104]) );
  XNOR2_X1 RoundFunction_T2_U258 ( .A(RoundFunction_STATE2[151]), .B(
        RoundFunction_T2_n572), .ZN(RoundFunction_TMP3_2[28]) );
  XNOR2_X1 RoundFunction_T2_U257 ( .A(RoundFunction_STATE2[150]), .B(
        RoundFunction_T2_n571), .ZN(RoundFunction_TMP3_2[27]) );
  XNOR2_X1 RoundFunction_T2_U256 ( .A(RoundFunction_STATE2[14]), .B(
        RoundFunction_T2_n594), .ZN(RoundFunction_TMP3_2[87]) );
  XNOR2_X1 RoundFunction_T2_U255 ( .A(RoundFunction_STATE2[149]), .B(
        RoundFunction_T2_n570), .ZN(RoundFunction_TMP3_2[26]) );
  XNOR2_X1 RoundFunction_T2_U254 ( .A(RoundFunction_STATE2[148]), .B(
        RoundFunction_T2_n569), .ZN(RoundFunction_TMP3_2[25]) );
  XNOR2_X1 RoundFunction_T2_U253 ( .A(RoundFunction_STATE2[147]), .B(
        RoundFunction_T2_n568), .ZN(RoundFunction_TMP3_2[24]) );
  XNOR2_X1 RoundFunction_T2_U252 ( .A(RoundFunction_STATE2[146]), .B(
        RoundFunction_T2_n567), .ZN(RoundFunction_TMP3_2[31]) );
  XNOR2_X1 RoundFunction_T2_U251 ( .A(RoundFunction_STATE2[145]), .B(
        RoundFunction_T2_n566), .ZN(RoundFunction_TMP3_2[30]) );
  XNOR2_X1 RoundFunction_T2_U250 ( .A(RoundFunction_STATE2[144]), .B(
        RoundFunction_T2_n565), .ZN(RoundFunction_TMP3_2[29]) );
  XNOR2_X1 RoundFunction_T2_U249 ( .A(RoundFunction_STATE2[143]), .B(
        RoundFunction_T2_n564), .ZN(RoundFunction_TMP3_2[150]) );
  XNOR2_X1 RoundFunction_T2_U248 ( .A(RoundFunction_STATE2[142]), .B(
        RoundFunction_T2_n563), .ZN(RoundFunction_TMP3_2[149]) );
  XNOR2_X1 RoundFunction_T2_U247 ( .A(RoundFunction_STATE2[141]), .B(
        RoundFunction_T2_n562), .ZN(RoundFunction_TMP3_2[148]) );
  XNOR2_X1 RoundFunction_T2_U246 ( .A(RoundFunction_STATE2[140]), .B(
        RoundFunction_T2_n561), .ZN(RoundFunction_TMP3_2[147]) );
  XNOR2_X1 RoundFunction_T2_U245 ( .A(RoundFunction_STATE2[13]), .B(
        RoundFunction_T2_n593), .ZN(RoundFunction_TMP3_2[86]) );
  XNOR2_X1 RoundFunction_T2_U244 ( .A(RoundFunction_STATE2[139]), .B(
        RoundFunction_T2_n599), .ZN(RoundFunction_TMP3_2[146]) );
  XNOR2_X1 RoundFunction_T2_U243 ( .A(RoundFunction_T2_n560), .B(
        RoundFunction_T2_n559), .ZN(RoundFunction_T2_n599) );
  XNOR2_X1 RoundFunction_T2_U242 ( .A(RoundFunction_STATE2[138]), .B(
        RoundFunction_T2_n598), .ZN(RoundFunction_TMP3_2[145]) );
  XNOR2_X1 RoundFunction_T2_U241 ( .A(RoundFunction_T2_n558), .B(
        RoundFunction_T2_n557), .ZN(RoundFunction_T2_n598) );
  XNOR2_X1 RoundFunction_T2_U240 ( .A(RoundFunction_STATE2[137]), .B(
        RoundFunction_T2_n597), .ZN(RoundFunction_TMP3_2[144]) );
  XNOR2_X1 RoundFunction_T2_U239 ( .A(RoundFunction_T2_n556), .B(
        RoundFunction_T2_n555), .ZN(RoundFunction_T2_n597) );
  XNOR2_X1 RoundFunction_T2_U238 ( .A(RoundFunction_STATE2[136]), .B(
        RoundFunction_T2_n596), .ZN(RoundFunction_TMP3_2[151]) );
  XNOR2_X1 RoundFunction_T2_U237 ( .A(RoundFunction_T2_n554), .B(
        RoundFunction_T2_n553), .ZN(RoundFunction_T2_n596) );
  XNOR2_X1 RoundFunction_T2_U236 ( .A(RoundFunction_STATE2[135]), .B(
        RoundFunction_T2_n595), .ZN(RoundFunction_TMP3_2[68]) );
  XNOR2_X1 RoundFunction_T2_U235 ( .A(RoundFunction_T2_n552), .B(
        RoundFunction_T2_n551), .ZN(RoundFunction_T2_n595) );
  XNOR2_X1 RoundFunction_T2_U234 ( .A(RoundFunction_STATE2[134]), .B(
        RoundFunction_T2_n594), .ZN(RoundFunction_TMP3_2[67]) );
  XNOR2_X1 RoundFunction_T2_U233 ( .A(RoundFunction_T2_n550), .B(
        RoundFunction_T2_n549), .ZN(RoundFunction_T2_n594) );
  XNOR2_X1 RoundFunction_T2_U232 ( .A(RoundFunction_STATE2[133]), .B(
        RoundFunction_T2_n593), .ZN(RoundFunction_TMP3_2[66]) );
  XNOR2_X1 RoundFunction_T2_U231 ( .A(RoundFunction_T2_n548), .B(
        RoundFunction_T2_n547), .ZN(RoundFunction_T2_n593) );
  XNOR2_X1 RoundFunction_T2_U230 ( .A(RoundFunction_STATE2[132]), .B(
        RoundFunction_T2_n592), .ZN(RoundFunction_TMP3_2[65]) );
  XNOR2_X1 RoundFunction_T2_U229 ( .A(RoundFunction_STATE2[131]), .B(
        RoundFunction_T2_n591), .ZN(RoundFunction_TMP3_2[64]) );
  XNOR2_X1 RoundFunction_T2_U228 ( .A(RoundFunction_STATE2[130]), .B(
        RoundFunction_T2_n590), .ZN(RoundFunction_TMP3_2[71]) );
  XNOR2_X1 RoundFunction_T2_U227 ( .A(RoundFunction_STATE2[12]), .B(
        RoundFunction_T2_n592), .ZN(RoundFunction_TMP3_2[85]) );
  XNOR2_X1 RoundFunction_T2_U226 ( .A(RoundFunction_T2_n546), .B(
        RoundFunction_T2_n545), .ZN(RoundFunction_T2_n592) );
  XNOR2_X1 RoundFunction_T2_U225 ( .A(RoundFunction_STATE2[129]), .B(
        RoundFunction_T2_n600), .ZN(RoundFunction_TMP3_2[70]) );
  XNOR2_X1 RoundFunction_T2_U224 ( .A(RoundFunction_T2_n544), .B(
        RoundFunction_T2_n543), .ZN(RoundFunction_T2_n600) );
  XNOR2_X1 RoundFunction_T2_U223 ( .A(RoundFunction_STATE2[128]), .B(
        RoundFunction_T2_n589), .ZN(RoundFunction_TMP3_2[69]) );
  XNOR2_X1 RoundFunction_T2_U222 ( .A(RoundFunction_T2_n542), .B(
        RoundFunction_T2_n541), .ZN(RoundFunction_T2_n589) );
  XNOR2_X1 RoundFunction_T2_U221 ( .A(RoundFunction_STATE2[127]), .B(
        RoundFunction_T2_n588), .ZN(RoundFunction_TMP3_2[184]) );
  XNOR2_X1 RoundFunction_T2_U220 ( .A(RoundFunction_T2_n540), .B(
        RoundFunction_T2_n539), .ZN(RoundFunction_T2_n588) );
  XNOR2_X1 RoundFunction_T2_U219 ( .A(RoundFunction_STATE2[126]), .B(
        RoundFunction_T2_n587), .ZN(RoundFunction_TMP3_2[191]) );
  XNOR2_X1 RoundFunction_T2_U218 ( .A(RoundFunction_T2_n538), .B(
        RoundFunction_T2_n537), .ZN(RoundFunction_T2_n587) );
  XNOR2_X1 RoundFunction_T2_U217 ( .A(RoundFunction_STATE2[125]), .B(
        RoundFunction_T2_n586), .ZN(RoundFunction_TMP3_2[190]) );
  XNOR2_X1 RoundFunction_T2_U216 ( .A(RoundFunction_T2_n536), .B(
        RoundFunction_T2_n535), .ZN(RoundFunction_T2_n586) );
  XNOR2_X1 RoundFunction_T2_U215 ( .A(RoundFunction_STATE2[124]), .B(
        RoundFunction_T2_n585), .ZN(RoundFunction_TMP3_2[189]) );
  XNOR2_X1 RoundFunction_T2_U214 ( .A(RoundFunction_T2_n534), .B(
        RoundFunction_T2_n559), .ZN(RoundFunction_T2_n585) );
  XOR2_X1 RoundFunction_T2_U213 ( .A(RoundFunction_STATE2[11]), .B(
        RoundFunction_T2_n533), .Z(RoundFunction_T2_n559) );
  XNOR2_X1 RoundFunction_T2_U212 ( .A(RoundFunction_T2_n532), .B(
        RoundFunction_T2_n531), .ZN(RoundFunction_T2_n533) );
  XNOR2_X1 RoundFunction_T2_U211 ( .A(RoundFunction_STATE2[51]), .B(
        RoundFunction_STATE2[91]), .ZN(RoundFunction_T2_n531) );
  XOR2_X1 RoundFunction_T2_U210 ( .A(RoundFunction_STATE2[131]), .B(
        RoundFunction_STATE2[171]), .Z(RoundFunction_T2_n532) );
  XNOR2_X1 RoundFunction_T2_U209 ( .A(RoundFunction_STATE2[123]), .B(
        RoundFunction_T2_n584), .ZN(RoundFunction_TMP3_2[188]) );
  XNOR2_X1 RoundFunction_T2_U208 ( .A(RoundFunction_T2_n530), .B(
        RoundFunction_T2_n557), .ZN(RoundFunction_T2_n584) );
  XOR2_X1 RoundFunction_T2_U207 ( .A(RoundFunction_STATE2[10]), .B(
        RoundFunction_T2_n529), .Z(RoundFunction_T2_n557) );
  XNOR2_X1 RoundFunction_T2_U206 ( .A(RoundFunction_T2_n528), .B(
        RoundFunction_T2_n527), .ZN(RoundFunction_T2_n529) );
  XNOR2_X1 RoundFunction_T2_U205 ( .A(RoundFunction_STATE2[50]), .B(
        RoundFunction_STATE2[90]), .ZN(RoundFunction_T2_n527) );
  XOR2_X1 RoundFunction_T2_U204 ( .A(RoundFunction_STATE2[130]), .B(
        RoundFunction_STATE2[170]), .Z(RoundFunction_T2_n528) );
  XNOR2_X1 RoundFunction_T2_U203 ( .A(RoundFunction_STATE2[122]), .B(
        RoundFunction_T2_n583), .ZN(RoundFunction_TMP3_2[187]) );
  XNOR2_X1 RoundFunction_T2_U202 ( .A(RoundFunction_T2_n526), .B(
        RoundFunction_T2_n555), .ZN(RoundFunction_T2_n583) );
  XOR2_X1 RoundFunction_T2_U201 ( .A(RoundFunction_STATE2[89]), .B(
        RoundFunction_T2_n525), .Z(RoundFunction_T2_n555) );
  XNOR2_X1 RoundFunction_T2_U200 ( .A(RoundFunction_T2_n524), .B(
        RoundFunction_T2_n523), .ZN(RoundFunction_T2_n525) );
  XNOR2_X1 RoundFunction_T2_U199 ( .A(RoundFunction_STATE2[129]), .B(
        RoundFunction_STATE2[49]), .ZN(RoundFunction_T2_n523) );
  XOR2_X1 RoundFunction_T2_U198 ( .A(RoundFunction_STATE2[169]), .B(
        RoundFunction_STATE2[9]), .Z(RoundFunction_T2_n524) );
  XNOR2_X1 RoundFunction_T2_U197 ( .A(RoundFunction_STATE2[121]), .B(
        RoundFunction_T2_n582), .ZN(RoundFunction_TMP3_2[186]) );
  XNOR2_X1 RoundFunction_T2_U196 ( .A(RoundFunction_T2_n522), .B(
        RoundFunction_T2_n553), .ZN(RoundFunction_T2_n582) );
  XOR2_X1 RoundFunction_T2_U195 ( .A(RoundFunction_STATE2[128]), .B(
        RoundFunction_T2_n521), .Z(RoundFunction_T2_n553) );
  XNOR2_X1 RoundFunction_T2_U194 ( .A(RoundFunction_T2_n520), .B(
        RoundFunction_T2_n519), .ZN(RoundFunction_T2_n521) );
  XNOR2_X1 RoundFunction_T2_U193 ( .A(RoundFunction_STATE2[48]), .B(
        RoundFunction_STATE2[8]), .ZN(RoundFunction_T2_n519) );
  XOR2_X1 RoundFunction_T2_U192 ( .A(RoundFunction_STATE2[88]), .B(
        RoundFunction_STATE2[168]), .Z(RoundFunction_T2_n520) );
  XNOR2_X1 RoundFunction_T2_U191 ( .A(RoundFunction_STATE2[120]), .B(
        RoundFunction_T2_n581), .ZN(RoundFunction_TMP3_2[185]) );
  XNOR2_X1 RoundFunction_T2_U190 ( .A(RoundFunction_STATE2[11]), .B(
        RoundFunction_T2_n591), .ZN(RoundFunction_TMP3_2[84]) );
  XNOR2_X1 RoundFunction_T2_U189 ( .A(RoundFunction_T2_n518), .B(
        RoundFunction_T2_n517), .ZN(RoundFunction_T2_n591) );
  XNOR2_X1 RoundFunction_T2_U188 ( .A(RoundFunction_STATE2[119]), .B(
        RoundFunction_T2_n580), .ZN(RoundFunction_TMP3_2[182]) );
  XNOR2_X1 RoundFunction_T2_U187 ( .A(RoundFunction_T2_n554), .B(
        RoundFunction_T2_n549), .ZN(RoundFunction_T2_n580) );
  XOR2_X1 RoundFunction_T2_U186 ( .A(RoundFunction_STATE2[126]), .B(
        RoundFunction_T2_n516), .Z(RoundFunction_T2_n549) );
  XNOR2_X1 RoundFunction_T2_U185 ( .A(RoundFunction_T2_n515), .B(
        RoundFunction_T2_n514), .ZN(RoundFunction_T2_n516) );
  XNOR2_X1 RoundFunction_T2_U184 ( .A(RoundFunction_STATE2[46]), .B(
        RoundFunction_STATE2[86]), .ZN(RoundFunction_T2_n514) );
  XOR2_X1 RoundFunction_T2_U183 ( .A(RoundFunction_STATE2[6]), .B(
        RoundFunction_STATE2[166]), .Z(RoundFunction_T2_n515) );
  XOR2_X1 RoundFunction_T2_U182 ( .A(RoundFunction_STATE2[111]), .B(
        RoundFunction_T2_n513), .Z(RoundFunction_T2_n554) );
  XNOR2_X1 RoundFunction_T2_U181 ( .A(RoundFunction_T2_n512), .B(
        RoundFunction_T2_n511), .ZN(RoundFunction_T2_n513) );
  XNOR2_X1 RoundFunction_T2_U180 ( .A(RoundFunction_STATE2[31]), .B(
        RoundFunction_STATE2[71]), .ZN(RoundFunction_T2_n511) );
  XOR2_X1 RoundFunction_T2_U179 ( .A(RoundFunction_STATE2[151]), .B(
        RoundFunction_STATE2[191]), .Z(RoundFunction_T2_n512) );
  XNOR2_X1 RoundFunction_T2_U178 ( .A(RoundFunction_STATE2[118]), .B(
        RoundFunction_T2_n579), .ZN(RoundFunction_TMP3_2[181]) );
  XNOR2_X1 RoundFunction_T2_U177 ( .A(RoundFunction_T2_n510), .B(
        RoundFunction_T2_n547), .ZN(RoundFunction_T2_n579) );
  XOR2_X1 RoundFunction_T2_U176 ( .A(RoundFunction_STATE2[125]), .B(
        RoundFunction_T2_n509), .Z(RoundFunction_T2_n547) );
  XNOR2_X1 RoundFunction_T2_U175 ( .A(RoundFunction_T2_n508), .B(
        RoundFunction_T2_n507), .ZN(RoundFunction_T2_n509) );
  XNOR2_X1 RoundFunction_T2_U174 ( .A(RoundFunction_STATE2[45]), .B(
        RoundFunction_STATE2[85]), .ZN(RoundFunction_T2_n507) );
  XOR2_X1 RoundFunction_T2_U173 ( .A(RoundFunction_STATE2[5]), .B(
        RoundFunction_STATE2[165]), .Z(RoundFunction_T2_n508) );
  XNOR2_X1 RoundFunction_T2_U172 ( .A(RoundFunction_STATE2[117]), .B(
        RoundFunction_T2_n578), .ZN(RoundFunction_TMP3_2[180]) );
  XNOR2_X1 RoundFunction_T2_U171 ( .A(RoundFunction_T2_n506), .B(
        RoundFunction_T2_n545), .ZN(RoundFunction_T2_n578) );
  XOR2_X1 RoundFunction_T2_U170 ( .A(RoundFunction_STATE2[124]), .B(
        RoundFunction_T2_n505), .Z(RoundFunction_T2_n545) );
  XNOR2_X1 RoundFunction_T2_U169 ( .A(RoundFunction_T2_n504), .B(
        RoundFunction_T2_n503), .ZN(RoundFunction_T2_n505) );
  XNOR2_X1 RoundFunction_T2_U168 ( .A(RoundFunction_STATE2[44]), .B(
        RoundFunction_STATE2[84]), .ZN(RoundFunction_T2_n503) );
  XOR2_X1 RoundFunction_T2_U167 ( .A(RoundFunction_STATE2[4]), .B(
        RoundFunction_STATE2[164]), .Z(RoundFunction_T2_n504) );
  XNOR2_X1 RoundFunction_T2_U166 ( .A(RoundFunction_STATE2[116]), .B(
        RoundFunction_T2_n577), .ZN(RoundFunction_TMP3_2[179]) );
  XNOR2_X1 RoundFunction_T2_U165 ( .A(RoundFunction_T2_n502), .B(
        RoundFunction_T2_n517), .ZN(RoundFunction_T2_n577) );
  XOR2_X1 RoundFunction_T2_U164 ( .A(RoundFunction_STATE2[123]), .B(
        RoundFunction_T2_n501), .Z(RoundFunction_T2_n517) );
  XNOR2_X1 RoundFunction_T2_U163 ( .A(RoundFunction_T2_n500), .B(
        RoundFunction_T2_n499), .ZN(RoundFunction_T2_n501) );
  XNOR2_X1 RoundFunction_T2_U162 ( .A(RoundFunction_STATE2[3]), .B(
        RoundFunction_STATE2[83]), .ZN(RoundFunction_T2_n499) );
  XOR2_X1 RoundFunction_T2_U161 ( .A(RoundFunction_STATE2[43]), .B(
        RoundFunction_STATE2[163]), .Z(RoundFunction_T2_n500) );
  XNOR2_X1 RoundFunction_T2_U160 ( .A(RoundFunction_STATE2[115]), .B(
        RoundFunction_T2_n576), .ZN(RoundFunction_TMP3_2[178]) );
  XNOR2_X1 RoundFunction_T2_U159 ( .A(RoundFunction_T2_n498), .B(
        RoundFunction_T2_n497), .ZN(RoundFunction_T2_n576) );
  XNOR2_X1 RoundFunction_T2_U158 ( .A(RoundFunction_STATE2[114]), .B(
        RoundFunction_T2_n575), .ZN(RoundFunction_TMP3_2[177]) );
  XNOR2_X1 RoundFunction_T2_U157 ( .A(RoundFunction_T2_n543), .B(
        RoundFunction_T2_n560), .ZN(RoundFunction_T2_n575) );
  XOR2_X1 RoundFunction_T2_U156 ( .A(RoundFunction_STATE2[106]), .B(
        RoundFunction_T2_n496), .Z(RoundFunction_T2_n560) );
  XNOR2_X1 RoundFunction_T2_U155 ( .A(RoundFunction_T2_n495), .B(
        RoundFunction_T2_n494), .ZN(RoundFunction_T2_n496) );
  XNOR2_X1 RoundFunction_T2_U154 ( .A(RoundFunction_STATE2[26]), .B(
        RoundFunction_STATE2[66]), .ZN(RoundFunction_T2_n494) );
  XOR2_X1 RoundFunction_T2_U153 ( .A(RoundFunction_STATE2[146]), .B(
        RoundFunction_STATE2[186]), .Z(RoundFunction_T2_n495) );
  XOR2_X1 RoundFunction_T2_U152 ( .A(RoundFunction_STATE2[121]), .B(
        RoundFunction_T2_n493), .Z(RoundFunction_T2_n543) );
  XNOR2_X1 RoundFunction_T2_U151 ( .A(RoundFunction_T2_n492), .B(
        RoundFunction_T2_n491), .ZN(RoundFunction_T2_n493) );
  XNOR2_X1 RoundFunction_T2_U150 ( .A(RoundFunction_STATE2[1]), .B(
        RoundFunction_STATE2[81]), .ZN(RoundFunction_T2_n491) );
  XOR2_X1 RoundFunction_T2_U149 ( .A(RoundFunction_STATE2[41]), .B(
        RoundFunction_STATE2[161]), .Z(RoundFunction_T2_n492) );
  XNOR2_X1 RoundFunction_T2_U148 ( .A(RoundFunction_STATE2[113]), .B(
        RoundFunction_T2_n574), .ZN(RoundFunction_TMP3_2[176]) );
  XNOR2_X1 RoundFunction_T2_U147 ( .A(RoundFunction_T2_n558), .B(
        RoundFunction_T2_n541), .ZN(RoundFunction_T2_n574) );
  XOR2_X1 RoundFunction_T2_U146 ( .A(RoundFunction_STATE2[0]), .B(
        RoundFunction_T2_n490), .Z(RoundFunction_T2_n541) );
  XNOR2_X1 RoundFunction_T2_U145 ( .A(RoundFunction_T2_n489), .B(
        RoundFunction_T2_n488), .ZN(RoundFunction_T2_n490) );
  XNOR2_X1 RoundFunction_T2_U144 ( .A(RoundFunction_STATE2[40]), .B(
        RoundFunction_STATE2[80]), .ZN(RoundFunction_T2_n488) );
  XOR2_X1 RoundFunction_T2_U143 ( .A(RoundFunction_STATE2[120]), .B(
        RoundFunction_STATE2[160]), .Z(RoundFunction_T2_n489) );
  XOR2_X1 RoundFunction_T2_U142 ( .A(RoundFunction_STATE2[105]), .B(
        RoundFunction_T2_n487), .Z(RoundFunction_T2_n558) );
  XNOR2_X1 RoundFunction_T2_U141 ( .A(RoundFunction_T2_n486), .B(
        RoundFunction_T2_n485), .ZN(RoundFunction_T2_n487) );
  XNOR2_X1 RoundFunction_T2_U140 ( .A(RoundFunction_STATE2[25]), .B(
        RoundFunction_STATE2[65]), .ZN(RoundFunction_T2_n485) );
  XOR2_X1 RoundFunction_T2_U139 ( .A(RoundFunction_STATE2[145]), .B(
        RoundFunction_STATE2[185]), .Z(RoundFunction_T2_n486) );
  XNOR2_X1 RoundFunction_T2_U138 ( .A(RoundFunction_STATE2[112]), .B(
        RoundFunction_T2_n573), .ZN(RoundFunction_TMP3_2[183]) );
  XNOR2_X1 RoundFunction_T2_U137 ( .A(RoundFunction_T2_n556), .B(
        RoundFunction_T2_n551), .ZN(RoundFunction_T2_n573) );
  XOR2_X1 RoundFunction_T2_U136 ( .A(RoundFunction_STATE2[127]), .B(
        RoundFunction_T2_n484), .Z(RoundFunction_T2_n551) );
  XNOR2_X1 RoundFunction_T2_U135 ( .A(RoundFunction_T2_n483), .B(
        RoundFunction_T2_n482), .ZN(RoundFunction_T2_n484) );
  XNOR2_X1 RoundFunction_T2_U134 ( .A(RoundFunction_STATE2[47]), .B(
        RoundFunction_STATE2[87]), .ZN(RoundFunction_T2_n482) );
  XOR2_X1 RoundFunction_T2_U133 ( .A(RoundFunction_STATE2[7]), .B(
        RoundFunction_STATE2[167]), .Z(RoundFunction_T2_n483) );
  XOR2_X1 RoundFunction_T2_U132 ( .A(RoundFunction_STATE2[104]), .B(
        RoundFunction_T2_n481), .Z(RoundFunction_T2_n556) );
  XNOR2_X1 RoundFunction_T2_U131 ( .A(RoundFunction_T2_n480), .B(
        RoundFunction_T2_n479), .ZN(RoundFunction_T2_n481) );
  XNOR2_X1 RoundFunction_T2_U130 ( .A(RoundFunction_STATE2[24]), .B(
        RoundFunction_STATE2[64]), .ZN(RoundFunction_T2_n479) );
  XOR2_X1 RoundFunction_T2_U129 ( .A(RoundFunction_STATE2[144]), .B(
        RoundFunction_STATE2[184]), .Z(RoundFunction_T2_n480) );
  XNOR2_X1 RoundFunction_T2_U128 ( .A(RoundFunction_STATE2[111]), .B(
        RoundFunction_T2_n572), .ZN(RoundFunction_TMP3_2[96]) );
  XNOR2_X1 RoundFunction_T2_U127 ( .A(RoundFunction_T2_n542), .B(
        RoundFunction_T2_n537), .ZN(RoundFunction_T2_n572) );
  XOR2_X1 RoundFunction_T2_U126 ( .A(RoundFunction_STATE2[118]), .B(
        RoundFunction_T2_n478), .Z(RoundFunction_T2_n537) );
  XNOR2_X1 RoundFunction_T2_U125 ( .A(RoundFunction_T2_n477), .B(
        RoundFunction_T2_n476), .ZN(RoundFunction_T2_n478) );
  XNOR2_X1 RoundFunction_T2_U124 ( .A(RoundFunction_STATE2[198]), .B(
        RoundFunction_STATE2[78]), .ZN(RoundFunction_T2_n476) );
  XOR2_X1 RoundFunction_T2_U123 ( .A(RoundFunction_STATE2[38]), .B(
        RoundFunction_STATE2[158]), .Z(RoundFunction_T2_n477) );
  XOR2_X1 RoundFunction_T2_U122 ( .A(RoundFunction_STATE2[103]), .B(
        RoundFunction_T2_n475), .Z(RoundFunction_T2_n542) );
  XNOR2_X1 RoundFunction_T2_U121 ( .A(RoundFunction_T2_n474), .B(
        RoundFunction_T2_n473), .ZN(RoundFunction_T2_n475) );
  XNOR2_X1 RoundFunction_T2_U120 ( .A(RoundFunction_STATE2[23]), .B(
        RoundFunction_STATE2[63]), .ZN(RoundFunction_T2_n473) );
  XOR2_X1 RoundFunction_T2_U119 ( .A(RoundFunction_STATE2[143]), .B(
        RoundFunction_STATE2[183]), .Z(RoundFunction_T2_n474) );
  XNOR2_X1 RoundFunction_T2_U118 ( .A(RoundFunction_STATE2[110]), .B(
        RoundFunction_T2_n571), .ZN(RoundFunction_TMP3_2[103]) );
  XNOR2_X1 RoundFunction_T2_U117 ( .A(RoundFunction_T2_n552), .B(
        RoundFunction_T2_n535), .ZN(RoundFunction_T2_n571) );
  XOR2_X1 RoundFunction_T2_U116 ( .A(RoundFunction_STATE2[117]), .B(
        RoundFunction_T2_n472), .Z(RoundFunction_T2_n535) );
  XNOR2_X1 RoundFunction_T2_U115 ( .A(RoundFunction_T2_n471), .B(
        RoundFunction_T2_n470), .ZN(RoundFunction_T2_n472) );
  XNOR2_X1 RoundFunction_T2_U114 ( .A(RoundFunction_STATE2[197]), .B(
        RoundFunction_STATE2[77]), .ZN(RoundFunction_T2_n470) );
  XOR2_X1 RoundFunction_T2_U113 ( .A(RoundFunction_STATE2[37]), .B(
        RoundFunction_STATE2[157]), .Z(RoundFunction_T2_n471) );
  XOR2_X1 RoundFunction_T2_U112 ( .A(RoundFunction_STATE2[102]), .B(
        RoundFunction_T2_n469), .Z(RoundFunction_T2_n552) );
  XNOR2_X1 RoundFunction_T2_U111 ( .A(RoundFunction_T2_n468), .B(
        RoundFunction_T2_n467), .ZN(RoundFunction_T2_n469) );
  XNOR2_X1 RoundFunction_T2_U110 ( .A(RoundFunction_STATE2[22]), .B(
        RoundFunction_STATE2[62]), .ZN(RoundFunction_T2_n467) );
  XOR2_X1 RoundFunction_T2_U109 ( .A(RoundFunction_STATE2[142]), .B(
        RoundFunction_STATE2[182]), .Z(RoundFunction_T2_n468) );
  XNOR2_X1 RoundFunction_T2_U108 ( .A(RoundFunction_STATE2[10]), .B(
        RoundFunction_T2_n590), .ZN(RoundFunction_TMP3_2[83]) );
  XNOR2_X1 RoundFunction_T2_U107 ( .A(RoundFunction_T2_n466), .B(
        RoundFunction_T2_n497), .ZN(RoundFunction_T2_n590) );
  XOR2_X1 RoundFunction_T2_U106 ( .A(RoundFunction_STATE2[122]), .B(
        RoundFunction_T2_n465), .Z(RoundFunction_T2_n497) );
  XNOR2_X1 RoundFunction_T2_U105 ( .A(RoundFunction_T2_n464), .B(
        RoundFunction_T2_n463), .ZN(RoundFunction_T2_n465) );
  XNOR2_X1 RoundFunction_T2_U104 ( .A(RoundFunction_STATE2[2]), .B(
        RoundFunction_STATE2[82]), .ZN(RoundFunction_T2_n463) );
  XOR2_X1 RoundFunction_T2_U103 ( .A(RoundFunction_STATE2[42]), .B(
        RoundFunction_STATE2[162]), .Z(RoundFunction_T2_n464) );
  XNOR2_X1 RoundFunction_T2_U102 ( .A(RoundFunction_STATE2[109]), .B(
        RoundFunction_T2_n570), .ZN(RoundFunction_TMP3_2[102]) );
  XNOR2_X1 RoundFunction_T2_U101 ( .A(RoundFunction_T2_n550), .B(
        RoundFunction_T2_n534), .ZN(RoundFunction_T2_n570) );
  XOR2_X1 RoundFunction_T2_U100 ( .A(RoundFunction_STATE2[116]), .B(
        RoundFunction_T2_n462), .Z(RoundFunction_T2_n534) );
  XNOR2_X1 RoundFunction_T2_U99 ( .A(RoundFunction_T2_n461), .B(
        RoundFunction_T2_n460), .ZN(RoundFunction_T2_n462) );
  XNOR2_X1 RoundFunction_T2_U98 ( .A(RoundFunction_STATE2[196]), .B(
        RoundFunction_STATE2[76]), .ZN(RoundFunction_T2_n460) );
  XOR2_X1 RoundFunction_T2_U97 ( .A(RoundFunction_STATE2[36]), .B(
        RoundFunction_STATE2[156]), .Z(RoundFunction_T2_n461) );
  XOR2_X1 RoundFunction_T2_U96 ( .A(RoundFunction_STATE2[101]), .B(
        RoundFunction_T2_n459), .Z(RoundFunction_T2_n550) );
  XNOR2_X1 RoundFunction_T2_U95 ( .A(RoundFunction_T2_n458), .B(
        RoundFunction_T2_n457), .ZN(RoundFunction_T2_n459) );
  XNOR2_X1 RoundFunction_T2_U94 ( .A(RoundFunction_STATE2[21]), .B(
        RoundFunction_STATE2[61]), .ZN(RoundFunction_T2_n457) );
  XOR2_X1 RoundFunction_T2_U93 ( .A(RoundFunction_STATE2[141]), .B(
        RoundFunction_STATE2[181]), .Z(RoundFunction_T2_n458) );
  XNOR2_X1 RoundFunction_T2_U92 ( .A(RoundFunction_STATE2[108]), .B(
        RoundFunction_T2_n569), .ZN(RoundFunction_TMP3_2[101]) );
  XNOR2_X1 RoundFunction_T2_U91 ( .A(RoundFunction_T2_n548), .B(
        RoundFunction_T2_n530), .ZN(RoundFunction_T2_n569) );
  XOR2_X1 RoundFunction_T2_U90 ( .A(RoundFunction_STATE2[115]), .B(
        RoundFunction_T2_n456), .Z(RoundFunction_T2_n530) );
  XNOR2_X1 RoundFunction_T2_U89 ( .A(RoundFunction_T2_n455), .B(
        RoundFunction_T2_n454), .ZN(RoundFunction_T2_n456) );
  XNOR2_X1 RoundFunction_T2_U88 ( .A(RoundFunction_STATE2[195]), .B(
        RoundFunction_STATE2[75]), .ZN(RoundFunction_T2_n454) );
  XOR2_X1 RoundFunction_T2_U87 ( .A(RoundFunction_STATE2[35]), .B(
        RoundFunction_STATE2[155]), .Z(RoundFunction_T2_n455) );
  XOR2_X1 RoundFunction_T2_U86 ( .A(RoundFunction_STATE2[100]), .B(
        RoundFunction_T2_n453), .Z(RoundFunction_T2_n548) );
  XNOR2_X1 RoundFunction_T2_U85 ( .A(RoundFunction_T2_n452), .B(
        RoundFunction_T2_n451), .ZN(RoundFunction_T2_n453) );
  XNOR2_X1 RoundFunction_T2_U84 ( .A(RoundFunction_STATE2[20]), .B(
        RoundFunction_STATE2[60]), .ZN(RoundFunction_T2_n451) );
  XOR2_X1 RoundFunction_T2_U83 ( .A(RoundFunction_STATE2[140]), .B(
        RoundFunction_STATE2[180]), .Z(RoundFunction_T2_n452) );
  XNOR2_X1 RoundFunction_T2_U82 ( .A(RoundFunction_STATE2[107]), .B(
        RoundFunction_T2_n568), .ZN(RoundFunction_TMP3_2[100]) );
  XNOR2_X1 RoundFunction_T2_U81 ( .A(RoundFunction_T2_n546), .B(
        RoundFunction_T2_n526), .ZN(RoundFunction_T2_n568) );
  XOR2_X1 RoundFunction_T2_U80 ( .A(RoundFunction_STATE2[114]), .B(
        RoundFunction_T2_n450), .Z(RoundFunction_T2_n526) );
  XNOR2_X1 RoundFunction_T2_U79 ( .A(RoundFunction_T2_n449), .B(
        RoundFunction_T2_n448), .ZN(RoundFunction_T2_n450) );
  XNOR2_X1 RoundFunction_T2_U78 ( .A(RoundFunction_STATE2[194]), .B(
        RoundFunction_STATE2[74]), .ZN(RoundFunction_T2_n448) );
  XOR2_X1 RoundFunction_T2_U77 ( .A(RoundFunction_STATE2[34]), .B(
        RoundFunction_STATE2[154]), .Z(RoundFunction_T2_n449) );
  XOR2_X1 RoundFunction_T2_U76 ( .A(RoundFunction_STATE2[59]), .B(
        RoundFunction_T2_n447), .Z(RoundFunction_T2_n546) );
  XNOR2_X1 RoundFunction_T2_U75 ( .A(RoundFunction_T2_n446), .B(
        RoundFunction_T2_n445), .ZN(RoundFunction_T2_n447) );
  XNOR2_X1 RoundFunction_T2_U74 ( .A(RoundFunction_STATE2[139]), .B(
        RoundFunction_STATE2[19]), .ZN(RoundFunction_T2_n445) );
  XOR2_X1 RoundFunction_T2_U73 ( .A(RoundFunction_STATE2[179]), .B(
        RoundFunction_STATE2[99]), .Z(RoundFunction_T2_n446) );
  XNOR2_X1 RoundFunction_T2_U72 ( .A(RoundFunction_STATE2[106]), .B(
        RoundFunction_T2_n567), .ZN(RoundFunction_TMP3_2[99]) );
  XNOR2_X1 RoundFunction_T2_U71 ( .A(RoundFunction_T2_n518), .B(
        RoundFunction_T2_n522), .ZN(RoundFunction_T2_n567) );
  XOR2_X1 RoundFunction_T2_U70 ( .A(RoundFunction_STATE2[113]), .B(
        RoundFunction_T2_n444), .Z(RoundFunction_T2_n522) );
  XNOR2_X1 RoundFunction_T2_U69 ( .A(RoundFunction_T2_n443), .B(
        RoundFunction_T2_n442), .ZN(RoundFunction_T2_n444) );
  XNOR2_X1 RoundFunction_T2_U68 ( .A(RoundFunction_STATE2[193]), .B(
        RoundFunction_STATE2[73]), .ZN(RoundFunction_T2_n442) );
  XOR2_X1 RoundFunction_T2_U67 ( .A(RoundFunction_STATE2[33]), .B(
        RoundFunction_STATE2[153]), .Z(RoundFunction_T2_n443) );
  XOR2_X1 RoundFunction_T2_U66 ( .A(RoundFunction_STATE2[58]), .B(
        RoundFunction_T2_n441), .Z(RoundFunction_T2_n518) );
  XNOR2_X1 RoundFunction_T2_U65 ( .A(RoundFunction_T2_n440), .B(
        RoundFunction_T2_n439), .ZN(RoundFunction_T2_n441) );
  XNOR2_X1 RoundFunction_T2_U64 ( .A(RoundFunction_STATE2[138]), .B(
        RoundFunction_STATE2[18]), .ZN(RoundFunction_T2_n439) );
  XOR2_X1 RoundFunction_T2_U63 ( .A(RoundFunction_STATE2[178]), .B(
        RoundFunction_STATE2[98]), .Z(RoundFunction_T2_n440) );
  XNOR2_X1 RoundFunction_T2_U62 ( .A(RoundFunction_STATE2[105]), .B(
        RoundFunction_T2_n566), .ZN(RoundFunction_TMP3_2[98]) );
  XNOR2_X1 RoundFunction_T2_U61 ( .A(RoundFunction_T2_n438), .B(
        RoundFunction_T2_n466), .ZN(RoundFunction_T2_n566) );
  XOR2_X1 RoundFunction_T2_U60 ( .A(RoundFunction_STATE2[57]), .B(
        RoundFunction_T2_n437), .Z(RoundFunction_T2_n466) );
  XNOR2_X1 RoundFunction_T2_U59 ( .A(RoundFunction_T2_n436), .B(
        RoundFunction_T2_n435), .ZN(RoundFunction_T2_n437) );
  XNOR2_X1 RoundFunction_T2_U58 ( .A(RoundFunction_STATE2[137]), .B(
        RoundFunction_STATE2[17]), .ZN(RoundFunction_T2_n435) );
  XOR2_X1 RoundFunction_T2_U57 ( .A(RoundFunction_STATE2[177]), .B(
        RoundFunction_STATE2[97]), .Z(RoundFunction_T2_n436) );
  XNOR2_X1 RoundFunction_T2_U56 ( .A(RoundFunction_STATE2[104]), .B(
        RoundFunction_T2_n565), .ZN(RoundFunction_TMP3_2[97]) );
  XNOR2_X1 RoundFunction_T2_U55 ( .A(RoundFunction_T2_n544), .B(
        RoundFunction_T2_n539), .ZN(RoundFunction_T2_n565) );
  XOR2_X1 RoundFunction_T2_U54 ( .A(RoundFunction_STATE2[119]), .B(
        RoundFunction_T2_n434), .Z(RoundFunction_T2_n539) );
  XNOR2_X1 RoundFunction_T2_U53 ( .A(RoundFunction_T2_n433), .B(
        RoundFunction_T2_n432), .ZN(RoundFunction_T2_n434) );
  XNOR2_X1 RoundFunction_T2_U52 ( .A(RoundFunction_STATE2[199]), .B(
        RoundFunction_STATE2[79]), .ZN(RoundFunction_T2_n432) );
  XOR2_X1 RoundFunction_T2_U51 ( .A(RoundFunction_STATE2[39]), .B(
        RoundFunction_STATE2[159]), .Z(RoundFunction_T2_n433) );
  XOR2_X1 RoundFunction_T2_U50 ( .A(RoundFunction_STATE2[136]), .B(
        RoundFunction_T2_n431), .Z(RoundFunction_T2_n544) );
  XNOR2_X1 RoundFunction_T2_U49 ( .A(RoundFunction_T2_n430), .B(
        RoundFunction_T2_n429), .ZN(RoundFunction_T2_n431) );
  XNOR2_X1 RoundFunction_T2_U48 ( .A(RoundFunction_STATE2[176]), .B(
        RoundFunction_STATE2[96]), .ZN(RoundFunction_T2_n429) );
  XOR2_X1 RoundFunction_T2_U47 ( .A(RoundFunction_STATE2[56]), .B(
        RoundFunction_STATE2[16]), .Z(RoundFunction_T2_n430) );
  XNOR2_X1 RoundFunction_T2_U46 ( .A(RoundFunction_STATE2[103]), .B(
        RoundFunction_T2_n564), .ZN(RoundFunction_TMP3_2[18]) );
  XNOR2_X1 RoundFunction_T2_U45 ( .A(RoundFunction_T2_n428), .B(
        RoundFunction_T2_n510), .ZN(RoundFunction_T2_n564) );
  XOR2_X1 RoundFunction_T2_U44 ( .A(RoundFunction_STATE2[110]), .B(
        RoundFunction_T2_n427), .Z(RoundFunction_T2_n510) );
  XNOR2_X1 RoundFunction_T2_U43 ( .A(RoundFunction_T2_n426), .B(
        RoundFunction_T2_n425), .ZN(RoundFunction_T2_n427) );
  XNOR2_X1 RoundFunction_T2_U42 ( .A(RoundFunction_STATE2[190]), .B(
        RoundFunction_STATE2[70]), .ZN(RoundFunction_T2_n425) );
  XOR2_X1 RoundFunction_T2_U41 ( .A(RoundFunction_STATE2[30]), .B(
        RoundFunction_STATE2[150]), .Z(RoundFunction_T2_n426) );
  XNOR2_X1 RoundFunction_T2_U40 ( .A(RoundFunction_STATE2[102]), .B(
        RoundFunction_T2_n563), .ZN(RoundFunction_TMP3_2[17]) );
  XNOR2_X1 RoundFunction_T2_U39 ( .A(RoundFunction_T2_n540), .B(
        RoundFunction_T2_n506), .ZN(RoundFunction_T2_n563) );
  XOR2_X1 RoundFunction_T2_U38 ( .A(RoundFunction_STATE2[109]), .B(
        RoundFunction_T2_n424), .Z(RoundFunction_T2_n506) );
  XNOR2_X1 RoundFunction_T2_U37 ( .A(RoundFunction_T2_n423), .B(
        RoundFunction_T2_n422), .ZN(RoundFunction_T2_n424) );
  XNOR2_X1 RoundFunction_T2_U36 ( .A(RoundFunction_STATE2[189]), .B(
        RoundFunction_STATE2[69]), .ZN(RoundFunction_T2_n422) );
  XOR2_X1 RoundFunction_T2_U35 ( .A(RoundFunction_STATE2[29]), .B(
        RoundFunction_STATE2[149]), .Z(RoundFunction_T2_n423) );
  XOR2_X1 RoundFunction_T2_U34 ( .A(RoundFunction_STATE2[54]), .B(
        RoundFunction_T2_n421), .Z(RoundFunction_T2_n540) );
  XNOR2_X1 RoundFunction_T2_U33 ( .A(RoundFunction_T2_n420), .B(
        RoundFunction_T2_n419), .ZN(RoundFunction_T2_n421) );
  XNOR2_X1 RoundFunction_T2_U32 ( .A(RoundFunction_STATE2[134]), .B(
        RoundFunction_STATE2[174]), .ZN(RoundFunction_T2_n419) );
  XOR2_X1 RoundFunction_T2_U31 ( .A(RoundFunction_STATE2[14]), .B(
        RoundFunction_STATE2[94]), .Z(RoundFunction_T2_n420) );
  XNOR2_X1 RoundFunction_T2_U30 ( .A(RoundFunction_STATE2[101]), .B(
        RoundFunction_T2_n562), .ZN(RoundFunction_TMP3_2[16]) );
  XNOR2_X1 RoundFunction_T2_U29 ( .A(RoundFunction_T2_n538), .B(
        RoundFunction_T2_n502), .ZN(RoundFunction_T2_n562) );
  XOR2_X1 RoundFunction_T2_U28 ( .A(RoundFunction_STATE2[108]), .B(
        RoundFunction_T2_n418), .Z(RoundFunction_T2_n502) );
  XNOR2_X1 RoundFunction_T2_U27 ( .A(RoundFunction_T2_n417), .B(
        RoundFunction_T2_n416), .ZN(RoundFunction_T2_n418) );
  XNOR2_X1 RoundFunction_T2_U26 ( .A(RoundFunction_STATE2[188]), .B(
        RoundFunction_STATE2[68]), .ZN(RoundFunction_T2_n416) );
  XOR2_X1 RoundFunction_T2_U25 ( .A(RoundFunction_STATE2[28]), .B(
        RoundFunction_STATE2[148]), .Z(RoundFunction_T2_n417) );
  XOR2_X1 RoundFunction_T2_U24 ( .A(RoundFunction_STATE2[53]), .B(
        RoundFunction_T2_n415), .Z(RoundFunction_T2_n538) );
  XNOR2_X1 RoundFunction_T2_U23 ( .A(RoundFunction_T2_n414), .B(
        RoundFunction_T2_n413), .ZN(RoundFunction_T2_n415) );
  XNOR2_X1 RoundFunction_T2_U22 ( .A(RoundFunction_STATE2[133]), .B(
        RoundFunction_STATE2[173]), .ZN(RoundFunction_T2_n413) );
  XOR2_X1 RoundFunction_T2_U21 ( .A(RoundFunction_STATE2[13]), .B(
        RoundFunction_STATE2[93]), .Z(RoundFunction_T2_n414) );
  XNOR2_X1 RoundFunction_T2_U20 ( .A(RoundFunction_STATE2[100]), .B(
        RoundFunction_T2_n561), .ZN(RoundFunction_TMP3_2[23]) );
  XNOR2_X1 RoundFunction_T2_U19 ( .A(RoundFunction_T2_n536), .B(
        RoundFunction_T2_n498), .ZN(RoundFunction_T2_n561) );
  XOR2_X1 RoundFunction_T2_U18 ( .A(RoundFunction_STATE2[107]), .B(
        RoundFunction_T2_n412), .Z(RoundFunction_T2_n498) );
  XNOR2_X1 RoundFunction_T2_U17 ( .A(RoundFunction_T2_n411), .B(
        RoundFunction_T2_n410), .ZN(RoundFunction_T2_n412) );
  XNOR2_X1 RoundFunction_T2_U16 ( .A(RoundFunction_STATE2[187]), .B(
        RoundFunction_STATE2[67]), .ZN(RoundFunction_T2_n410) );
  XOR2_X1 RoundFunction_T2_U15 ( .A(RoundFunction_STATE2[27]), .B(
        RoundFunction_STATE2[147]), .Z(RoundFunction_T2_n411) );
  XOR2_X1 RoundFunction_T2_U14 ( .A(RoundFunction_STATE2[52]), .B(
        RoundFunction_T2_n409), .Z(RoundFunction_T2_n536) );
  XNOR2_X1 RoundFunction_T2_U13 ( .A(RoundFunction_T2_n408), .B(
        RoundFunction_T2_n407), .ZN(RoundFunction_T2_n409) );
  XNOR2_X1 RoundFunction_T2_U12 ( .A(RoundFunction_STATE2[12]), .B(
        RoundFunction_STATE2[172]), .ZN(RoundFunction_T2_n407) );
  XOR2_X1 RoundFunction_T2_U11 ( .A(RoundFunction_STATE2[132]), .B(
        RoundFunction_STATE2[92]), .Z(RoundFunction_T2_n408) );
  XNOR2_X1 RoundFunction_T2_U10 ( .A(RoundFunction_STATE2[0]), .B(
        RoundFunction_T2_n581), .ZN(RoundFunction_TMP3_2[0]) );
  XNOR2_X1 RoundFunction_T2_U9 ( .A(RoundFunction_T2_n438), .B(
        RoundFunction_T2_n428), .ZN(RoundFunction_T2_n581) );
  XOR2_X1 RoundFunction_T2_U8 ( .A(RoundFunction_STATE2[55]), .B(
        RoundFunction_T2_n406), .Z(RoundFunction_T2_n428) );
  XNOR2_X1 RoundFunction_T2_U7 ( .A(RoundFunction_T2_n405), .B(
        RoundFunction_T2_n404), .ZN(RoundFunction_T2_n406) );
  XNOR2_X1 RoundFunction_T2_U6 ( .A(RoundFunction_STATE2[135]), .B(
        RoundFunction_STATE2[175]), .ZN(RoundFunction_T2_n404) );
  XOR2_X1 RoundFunction_T2_U5 ( .A(RoundFunction_STATE2[15]), .B(
        RoundFunction_STATE2[95]), .Z(RoundFunction_T2_n405) );
  XOR2_X1 RoundFunction_T2_U4 ( .A(RoundFunction_STATE2[112]), .B(
        RoundFunction_T2_n403), .Z(RoundFunction_T2_n438) );
  XNOR2_X1 RoundFunction_T2_U3 ( .A(RoundFunction_T2_n402), .B(
        RoundFunction_T2_n401), .ZN(RoundFunction_T2_n403) );
  XNOR2_X1 RoundFunction_T2_U2 ( .A(RoundFunction_STATE2[192]), .B(
        RoundFunction_STATE2[72]), .ZN(RoundFunction_T2_n401) );
  XOR2_X1 RoundFunction_T2_U1 ( .A(RoundFunction_STATE2[32]), .B(
        RoundFunction_STATE2[152]), .Z(RoundFunction_T2_n402) );
  XNOR2_X1 RoundFunction_T3_U400 ( .A(RoundFunction_STATE3[9]), .B(
        RoundFunction_T3_n600), .ZN(RoundFunction_TMP3_3[82]) );
  XNOR2_X1 RoundFunction_T3_U399 ( .A(RoundFunction_STATE3[99]), .B(
        RoundFunction_T3_n599), .ZN(RoundFunction_TMP3_3[22]) );
  XNOR2_X1 RoundFunction_T3_U398 ( .A(RoundFunction_STATE3[98]), .B(
        RoundFunction_T3_n598), .ZN(RoundFunction_TMP3_3[21]) );
  XNOR2_X1 RoundFunction_T3_U397 ( .A(RoundFunction_STATE3[97]), .B(
        RoundFunction_T3_n597), .ZN(RoundFunction_TMP3_3[20]) );
  XNOR2_X1 RoundFunction_T3_U396 ( .A(RoundFunction_STATE3[96]), .B(
        RoundFunction_T3_n596), .ZN(RoundFunction_TMP3_3[19]) );
  XNOR2_X1 RoundFunction_T3_U395 ( .A(RoundFunction_STATE3[95]), .B(
        RoundFunction_T3_n595), .ZN(RoundFunction_TMP3_3[137]) );
  XNOR2_X1 RoundFunction_T3_U394 ( .A(RoundFunction_STATE3[94]), .B(
        RoundFunction_T3_n594), .ZN(RoundFunction_TMP3_3[136]) );
  XNOR2_X1 RoundFunction_T3_U393 ( .A(RoundFunction_STATE3[93]), .B(
        RoundFunction_T3_n593), .ZN(RoundFunction_TMP3_3[143]) );
  XNOR2_X1 RoundFunction_T3_U392 ( .A(RoundFunction_STATE3[92]), .B(
        RoundFunction_T3_n592), .ZN(RoundFunction_TMP3_3[142]) );
  XNOR2_X1 RoundFunction_T3_U391 ( .A(RoundFunction_STATE3[91]), .B(
        RoundFunction_T3_n591), .ZN(RoundFunction_TMP3_3[141]) );
  XNOR2_X1 RoundFunction_T3_U390 ( .A(RoundFunction_STATE3[90]), .B(
        RoundFunction_T3_n590), .ZN(RoundFunction_TMP3_3[140]) );
  XNOR2_X1 RoundFunction_T3_U389 ( .A(RoundFunction_STATE3[8]), .B(
        RoundFunction_T3_n589), .ZN(RoundFunction_TMP3_3[81]) );
  XNOR2_X1 RoundFunction_T3_U388 ( .A(RoundFunction_STATE3[89]), .B(
        RoundFunction_T3_n600), .ZN(RoundFunction_TMP3_3[139]) );
  XNOR2_X1 RoundFunction_T3_U387 ( .A(RoundFunction_STATE3[88]), .B(
        RoundFunction_T3_n589), .ZN(RoundFunction_TMP3_3[138]) );
  XNOR2_X1 RoundFunction_T3_U386 ( .A(RoundFunction_STATE3[87]), .B(
        RoundFunction_T3_n588), .ZN(RoundFunction_TMP3_3[58]) );
  XNOR2_X1 RoundFunction_T3_U385 ( .A(RoundFunction_STATE3[86]), .B(
        RoundFunction_T3_n587), .ZN(RoundFunction_TMP3_3[57]) );
  XNOR2_X1 RoundFunction_T3_U384 ( .A(RoundFunction_STATE3[85]), .B(
        RoundFunction_T3_n586), .ZN(RoundFunction_TMP3_3[56]) );
  XNOR2_X1 RoundFunction_T3_U383 ( .A(RoundFunction_STATE3[84]), .B(
        RoundFunction_T3_n585), .ZN(RoundFunction_TMP3_3[63]) );
  XNOR2_X1 RoundFunction_T3_U382 ( .A(RoundFunction_STATE3[83]), .B(
        RoundFunction_T3_n584), .ZN(RoundFunction_TMP3_3[62]) );
  XNOR2_X1 RoundFunction_T3_U381 ( .A(RoundFunction_STATE3[82]), .B(
        RoundFunction_T3_n583), .ZN(RoundFunction_TMP3_3[61]) );
  XNOR2_X1 RoundFunction_T3_U380 ( .A(RoundFunction_STATE3[81]), .B(
        RoundFunction_T3_n582), .ZN(RoundFunction_TMP3_3[60]) );
  XNOR2_X1 RoundFunction_T3_U379 ( .A(RoundFunction_STATE3[80]), .B(
        RoundFunction_T3_n581), .ZN(RoundFunction_TMP3_3[59]) );
  XNOR2_X1 RoundFunction_T3_U378 ( .A(RoundFunction_STATE3[7]), .B(
        RoundFunction_T3_n588), .ZN(RoundFunction_TMP3_3[7]) );
  XNOR2_X1 RoundFunction_T3_U377 ( .A(RoundFunction_STATE3[79]), .B(
        RoundFunction_T3_n580), .ZN(RoundFunction_TMP3_3[51]) );
  XNOR2_X1 RoundFunction_T3_U376 ( .A(RoundFunction_STATE3[78]), .B(
        RoundFunction_T3_n579), .ZN(RoundFunction_TMP3_3[50]) );
  XNOR2_X1 RoundFunction_T3_U375 ( .A(RoundFunction_STATE3[77]), .B(
        RoundFunction_T3_n578), .ZN(RoundFunction_TMP3_3[49]) );
  XNOR2_X1 RoundFunction_T3_U374 ( .A(RoundFunction_STATE3[76]), .B(
        RoundFunction_T3_n577), .ZN(RoundFunction_TMP3_3[48]) );
  XNOR2_X1 RoundFunction_T3_U373 ( .A(RoundFunction_STATE3[75]), .B(
        RoundFunction_T3_n576), .ZN(RoundFunction_TMP3_3[55]) );
  XNOR2_X1 RoundFunction_T3_U372 ( .A(RoundFunction_STATE3[74]), .B(
        RoundFunction_T3_n575), .ZN(RoundFunction_TMP3_3[54]) );
  XNOR2_X1 RoundFunction_T3_U371 ( .A(RoundFunction_STATE3[73]), .B(
        RoundFunction_T3_n574), .ZN(RoundFunction_TMP3_3[53]) );
  XNOR2_X1 RoundFunction_T3_U370 ( .A(RoundFunction_STATE3[72]), .B(
        RoundFunction_T3_n573), .ZN(RoundFunction_TMP3_3[52]) );
  XNOR2_X1 RoundFunction_T3_U369 ( .A(RoundFunction_STATE3[71]), .B(
        RoundFunction_T3_n572), .ZN(RoundFunction_TMP3_3[174]) );
  XNOR2_X1 RoundFunction_T3_U368 ( .A(RoundFunction_STATE3[70]), .B(
        RoundFunction_T3_n571), .ZN(RoundFunction_TMP3_3[173]) );
  XNOR2_X1 RoundFunction_T3_U367 ( .A(RoundFunction_STATE3[6]), .B(
        RoundFunction_T3_n587), .ZN(RoundFunction_TMP3_3[6]) );
  XNOR2_X1 RoundFunction_T3_U366 ( .A(RoundFunction_STATE3[69]), .B(
        RoundFunction_T3_n570), .ZN(RoundFunction_TMP3_3[172]) );
  XNOR2_X1 RoundFunction_T3_U365 ( .A(RoundFunction_STATE3[68]), .B(
        RoundFunction_T3_n569), .ZN(RoundFunction_TMP3_3[171]) );
  XNOR2_X1 RoundFunction_T3_U364 ( .A(RoundFunction_STATE3[67]), .B(
        RoundFunction_T3_n568), .ZN(RoundFunction_TMP3_3[170]) );
  XNOR2_X1 RoundFunction_T3_U363 ( .A(RoundFunction_STATE3[66]), .B(
        RoundFunction_T3_n567), .ZN(RoundFunction_TMP3_3[169]) );
  XNOR2_X1 RoundFunction_T3_U362 ( .A(RoundFunction_STATE3[65]), .B(
        RoundFunction_T3_n566), .ZN(RoundFunction_TMP3_3[168]) );
  XNOR2_X1 RoundFunction_T3_U361 ( .A(RoundFunction_STATE3[64]), .B(
        RoundFunction_T3_n565), .ZN(RoundFunction_TMP3_3[175]) );
  XNOR2_X1 RoundFunction_T3_U360 ( .A(RoundFunction_STATE3[63]), .B(
        RoundFunction_T3_n564), .ZN(RoundFunction_TMP3_3[93]) );
  XNOR2_X1 RoundFunction_T3_U359 ( .A(RoundFunction_STATE3[62]), .B(
        RoundFunction_T3_n563), .ZN(RoundFunction_TMP3_3[92]) );
  XNOR2_X1 RoundFunction_T3_U358 ( .A(RoundFunction_STATE3[61]), .B(
        RoundFunction_T3_n562), .ZN(RoundFunction_TMP3_3[91]) );
  XNOR2_X1 RoundFunction_T3_U357 ( .A(RoundFunction_STATE3[60]), .B(
        RoundFunction_T3_n561), .ZN(RoundFunction_TMP3_3[90]) );
  XNOR2_X1 RoundFunction_T3_U356 ( .A(RoundFunction_STATE3[5]), .B(
        RoundFunction_T3_n586), .ZN(RoundFunction_TMP3_3[5]) );
  XNOR2_X1 RoundFunction_T3_U355 ( .A(RoundFunction_STATE3[59]), .B(
        RoundFunction_T3_n599), .ZN(RoundFunction_TMP3_3[89]) );
  XNOR2_X1 RoundFunction_T3_U354 ( .A(RoundFunction_STATE3[58]), .B(
        RoundFunction_T3_n598), .ZN(RoundFunction_TMP3_3[88]) );
  XNOR2_X1 RoundFunction_T3_U353 ( .A(RoundFunction_STATE3[57]), .B(
        RoundFunction_T3_n597), .ZN(RoundFunction_TMP3_3[95]) );
  XNOR2_X1 RoundFunction_T3_U352 ( .A(RoundFunction_STATE3[56]), .B(
        RoundFunction_T3_n596), .ZN(RoundFunction_TMP3_3[94]) );
  XNOR2_X1 RoundFunction_T3_U351 ( .A(RoundFunction_STATE3[55]), .B(
        RoundFunction_T3_n595), .ZN(RoundFunction_TMP3_3[11]) );
  XNOR2_X1 RoundFunction_T3_U350 ( .A(RoundFunction_STATE3[54]), .B(
        RoundFunction_T3_n594), .ZN(RoundFunction_TMP3_3[10]) );
  XNOR2_X1 RoundFunction_T3_U349 ( .A(RoundFunction_STATE3[53]), .B(
        RoundFunction_T3_n593), .ZN(RoundFunction_TMP3_3[9]) );
  XNOR2_X1 RoundFunction_T3_U348 ( .A(RoundFunction_STATE3[52]), .B(
        RoundFunction_T3_n592), .ZN(RoundFunction_TMP3_3[8]) );
  XNOR2_X1 RoundFunction_T3_U347 ( .A(RoundFunction_STATE3[51]), .B(
        RoundFunction_T3_n591), .ZN(RoundFunction_TMP3_3[15]) );
  XNOR2_X1 RoundFunction_T3_U346 ( .A(RoundFunction_STATE3[50]), .B(
        RoundFunction_T3_n590), .ZN(RoundFunction_TMP3_3[14]) );
  XNOR2_X1 RoundFunction_T3_U345 ( .A(RoundFunction_STATE3[4]), .B(
        RoundFunction_T3_n585), .ZN(RoundFunction_TMP3_3[4]) );
  XNOR2_X1 RoundFunction_T3_U344 ( .A(RoundFunction_STATE3[49]), .B(
        RoundFunction_T3_n600), .ZN(RoundFunction_TMP3_3[13]) );
  XNOR2_X1 RoundFunction_T3_U343 ( .A(RoundFunction_STATE3[48]), .B(
        RoundFunction_T3_n589), .ZN(RoundFunction_TMP3_3[12]) );
  XNOR2_X1 RoundFunction_T3_U342 ( .A(RoundFunction_STATE3[47]), .B(
        RoundFunction_T3_n588), .ZN(RoundFunction_TMP3_3[131]) );
  XNOR2_X1 RoundFunction_T3_U341 ( .A(RoundFunction_STATE3[46]), .B(
        RoundFunction_T3_n587), .ZN(RoundFunction_TMP3_3[130]) );
  XNOR2_X1 RoundFunction_T3_U340 ( .A(RoundFunction_STATE3[45]), .B(
        RoundFunction_T3_n586), .ZN(RoundFunction_TMP3_3[129]) );
  XNOR2_X1 RoundFunction_T3_U339 ( .A(RoundFunction_STATE3[44]), .B(
        RoundFunction_T3_n585), .ZN(RoundFunction_TMP3_3[128]) );
  XNOR2_X1 RoundFunction_T3_U338 ( .A(RoundFunction_STATE3[43]), .B(
        RoundFunction_T3_n584), .ZN(RoundFunction_TMP3_3[135]) );
  XNOR2_X1 RoundFunction_T3_U337 ( .A(RoundFunction_STATE3[42]), .B(
        RoundFunction_T3_n583), .ZN(RoundFunction_TMP3_3[134]) );
  XNOR2_X1 RoundFunction_T3_U336 ( .A(RoundFunction_STATE3[41]), .B(
        RoundFunction_T3_n582), .ZN(RoundFunction_TMP3_3[133]) );
  XNOR2_X1 RoundFunction_T3_U335 ( .A(RoundFunction_STATE3[40]), .B(
        RoundFunction_T3_n581), .ZN(RoundFunction_TMP3_3[132]) );
  XNOR2_X1 RoundFunction_T3_U334 ( .A(RoundFunction_STATE3[3]), .B(
        RoundFunction_T3_n584), .ZN(RoundFunction_TMP3_3[3]) );
  XNOR2_X1 RoundFunction_T3_U333 ( .A(RoundFunction_STATE3[39]), .B(
        RoundFunction_T3_n580), .ZN(RoundFunction_TMP3_3[122]) );
  XNOR2_X1 RoundFunction_T3_U332 ( .A(RoundFunction_STATE3[38]), .B(
        RoundFunction_T3_n579), .ZN(RoundFunction_TMP3_3[121]) );
  XNOR2_X1 RoundFunction_T3_U331 ( .A(RoundFunction_STATE3[37]), .B(
        RoundFunction_T3_n578), .ZN(RoundFunction_TMP3_3[120]) );
  XNOR2_X1 RoundFunction_T3_U330 ( .A(RoundFunction_STATE3[36]), .B(
        RoundFunction_T3_n577), .ZN(RoundFunction_TMP3_3[127]) );
  XNOR2_X1 RoundFunction_T3_U329 ( .A(RoundFunction_STATE3[35]), .B(
        RoundFunction_T3_n576), .ZN(RoundFunction_TMP3_3[126]) );
  XNOR2_X1 RoundFunction_T3_U328 ( .A(RoundFunction_STATE3[34]), .B(
        RoundFunction_T3_n575), .ZN(RoundFunction_TMP3_3[125]) );
  XNOR2_X1 RoundFunction_T3_U327 ( .A(RoundFunction_STATE3[33]), .B(
        RoundFunction_T3_n574), .ZN(RoundFunction_TMP3_3[124]) );
  XNOR2_X1 RoundFunction_T3_U326 ( .A(RoundFunction_STATE3[32]), .B(
        RoundFunction_T3_n573), .ZN(RoundFunction_TMP3_3[123]) );
  XNOR2_X1 RoundFunction_T3_U325 ( .A(RoundFunction_STATE3[31]), .B(
        RoundFunction_T3_n572), .ZN(RoundFunction_TMP3_3[43]) );
  XNOR2_X1 RoundFunction_T3_U324 ( .A(RoundFunction_STATE3[30]), .B(
        RoundFunction_T3_n571), .ZN(RoundFunction_TMP3_3[42]) );
  XNOR2_X1 RoundFunction_T3_U323 ( .A(RoundFunction_STATE3[2]), .B(
        RoundFunction_T3_n583), .ZN(RoundFunction_TMP3_3[2]) );
  XNOR2_X1 RoundFunction_T3_U322 ( .A(RoundFunction_STATE3[29]), .B(
        RoundFunction_T3_n570), .ZN(RoundFunction_TMP3_3[41]) );
  XNOR2_X1 RoundFunction_T3_U321 ( .A(RoundFunction_STATE3[28]), .B(
        RoundFunction_T3_n569), .ZN(RoundFunction_TMP3_3[40]) );
  XNOR2_X1 RoundFunction_T3_U320 ( .A(RoundFunction_STATE3[27]), .B(
        RoundFunction_T3_n568), .ZN(RoundFunction_TMP3_3[47]) );
  XNOR2_X1 RoundFunction_T3_U319 ( .A(RoundFunction_STATE3[26]), .B(
        RoundFunction_T3_n567), .ZN(RoundFunction_TMP3_3[46]) );
  XNOR2_X1 RoundFunction_T3_U318 ( .A(RoundFunction_STATE3[25]), .B(
        RoundFunction_T3_n566), .ZN(RoundFunction_TMP3_3[45]) );
  XNOR2_X1 RoundFunction_T3_U317 ( .A(RoundFunction_STATE3[24]), .B(
        RoundFunction_T3_n565), .ZN(RoundFunction_TMP3_3[44]) );
  XNOR2_X1 RoundFunction_T3_U316 ( .A(RoundFunction_STATE3[23]), .B(
        RoundFunction_T3_n564), .ZN(RoundFunction_TMP3_3[165]) );
  XNOR2_X1 RoundFunction_T3_U315 ( .A(RoundFunction_STATE3[22]), .B(
        RoundFunction_T3_n563), .ZN(RoundFunction_TMP3_3[164]) );
  XNOR2_X1 RoundFunction_T3_U314 ( .A(RoundFunction_STATE3[21]), .B(
        RoundFunction_T3_n562), .ZN(RoundFunction_TMP3_3[163]) );
  XNOR2_X1 RoundFunction_T3_U313 ( .A(RoundFunction_STATE3[20]), .B(
        RoundFunction_T3_n561), .ZN(RoundFunction_TMP3_3[162]) );
  XNOR2_X1 RoundFunction_T3_U312 ( .A(RoundFunction_STATE3[1]), .B(
        RoundFunction_T3_n582), .ZN(RoundFunction_TMP3_3[1]) );
  XNOR2_X1 RoundFunction_T3_U311 ( .A(RoundFunction_STATE3[19]), .B(
        RoundFunction_T3_n599), .ZN(RoundFunction_TMP3_3[161]) );
  XNOR2_X1 RoundFunction_T3_U310 ( .A(RoundFunction_STATE3[199]), .B(
        RoundFunction_T3_n580), .ZN(RoundFunction_TMP3_3[37]) );
  XNOR2_X1 RoundFunction_T3_U309 ( .A(RoundFunction_STATE3[198]), .B(
        RoundFunction_T3_n579), .ZN(RoundFunction_TMP3_3[36]) );
  XNOR2_X1 RoundFunction_T3_U308 ( .A(RoundFunction_STATE3[197]), .B(
        RoundFunction_T3_n578), .ZN(RoundFunction_TMP3_3[35]) );
  XNOR2_X1 RoundFunction_T3_U307 ( .A(RoundFunction_STATE3[196]), .B(
        RoundFunction_T3_n577), .ZN(RoundFunction_TMP3_3[34]) );
  XNOR2_X1 RoundFunction_T3_U306 ( .A(RoundFunction_STATE3[195]), .B(
        RoundFunction_T3_n576), .ZN(RoundFunction_TMP3_3[33]) );
  XNOR2_X1 RoundFunction_T3_U305 ( .A(RoundFunction_STATE3[194]), .B(
        RoundFunction_T3_n575), .ZN(RoundFunction_TMP3_3[32]) );
  XNOR2_X1 RoundFunction_T3_U304 ( .A(RoundFunction_STATE3[193]), .B(
        RoundFunction_T3_n574), .ZN(RoundFunction_TMP3_3[39]) );
  XNOR2_X1 RoundFunction_T3_U303 ( .A(RoundFunction_STATE3[192]), .B(
        RoundFunction_T3_n573), .ZN(RoundFunction_TMP3_3[38]) );
  XNOR2_X1 RoundFunction_T3_U302 ( .A(RoundFunction_STATE3[191]), .B(
        RoundFunction_T3_n572), .ZN(RoundFunction_TMP3_3[159]) );
  XNOR2_X1 RoundFunction_T3_U301 ( .A(RoundFunction_STATE3[190]), .B(
        RoundFunction_T3_n571), .ZN(RoundFunction_TMP3_3[158]) );
  XNOR2_X1 RoundFunction_T3_U300 ( .A(RoundFunction_STATE3[18]), .B(
        RoundFunction_T3_n598), .ZN(RoundFunction_TMP3_3[160]) );
  XNOR2_X1 RoundFunction_T3_U299 ( .A(RoundFunction_STATE3[189]), .B(
        RoundFunction_T3_n570), .ZN(RoundFunction_TMP3_3[157]) );
  XNOR2_X1 RoundFunction_T3_U298 ( .A(RoundFunction_STATE3[188]), .B(
        RoundFunction_T3_n569), .ZN(RoundFunction_TMP3_3[156]) );
  XNOR2_X1 RoundFunction_T3_U297 ( .A(RoundFunction_STATE3[187]), .B(
        RoundFunction_T3_n568), .ZN(RoundFunction_TMP3_3[155]) );
  XNOR2_X1 RoundFunction_T3_U296 ( .A(RoundFunction_STATE3[186]), .B(
        RoundFunction_T3_n567), .ZN(RoundFunction_TMP3_3[154]) );
  XNOR2_X1 RoundFunction_T3_U295 ( .A(RoundFunction_STATE3[185]), .B(
        RoundFunction_T3_n566), .ZN(RoundFunction_TMP3_3[153]) );
  XNOR2_X1 RoundFunction_T3_U294 ( .A(RoundFunction_STATE3[184]), .B(
        RoundFunction_T3_n565), .ZN(RoundFunction_TMP3_3[152]) );
  XNOR2_X1 RoundFunction_T3_U293 ( .A(RoundFunction_STATE3[183]), .B(
        RoundFunction_T3_n564), .ZN(RoundFunction_TMP3_3[76]) );
  XNOR2_X1 RoundFunction_T3_U292 ( .A(RoundFunction_STATE3[182]), .B(
        RoundFunction_T3_n563), .ZN(RoundFunction_TMP3_3[75]) );
  XNOR2_X1 RoundFunction_T3_U291 ( .A(RoundFunction_STATE3[181]), .B(
        RoundFunction_T3_n562), .ZN(RoundFunction_TMP3_3[74]) );
  XNOR2_X1 RoundFunction_T3_U290 ( .A(RoundFunction_STATE3[180]), .B(
        RoundFunction_T3_n561), .ZN(RoundFunction_TMP3_3[73]) );
  XNOR2_X1 RoundFunction_T3_U289 ( .A(RoundFunction_STATE3[17]), .B(
        RoundFunction_T3_n597), .ZN(RoundFunction_TMP3_3[167]) );
  XNOR2_X1 RoundFunction_T3_U288 ( .A(RoundFunction_STATE3[179]), .B(
        RoundFunction_T3_n599), .ZN(RoundFunction_TMP3_3[72]) );
  XNOR2_X1 RoundFunction_T3_U287 ( .A(RoundFunction_STATE3[178]), .B(
        RoundFunction_T3_n598), .ZN(RoundFunction_TMP3_3[79]) );
  XNOR2_X1 RoundFunction_T3_U286 ( .A(RoundFunction_STATE3[177]), .B(
        RoundFunction_T3_n597), .ZN(RoundFunction_TMP3_3[78]) );
  XNOR2_X1 RoundFunction_T3_U285 ( .A(RoundFunction_STATE3[176]), .B(
        RoundFunction_T3_n596), .ZN(RoundFunction_TMP3_3[77]) );
  XNOR2_X1 RoundFunction_T3_U284 ( .A(RoundFunction_STATE3[175]), .B(
        RoundFunction_T3_n595), .ZN(RoundFunction_TMP3_3[193]) );
  XNOR2_X1 RoundFunction_T3_U283 ( .A(RoundFunction_STATE3[174]), .B(
        RoundFunction_T3_n594), .ZN(RoundFunction_TMP3_3[192]) );
  XNOR2_X1 RoundFunction_T3_U282 ( .A(RoundFunction_STATE3[173]), .B(
        RoundFunction_T3_n593), .ZN(RoundFunction_TMP3_3[199]) );
  XNOR2_X1 RoundFunction_T3_U281 ( .A(RoundFunction_STATE3[172]), .B(
        RoundFunction_T3_n592), .ZN(RoundFunction_TMP3_3[198]) );
  XNOR2_X1 RoundFunction_T3_U280 ( .A(RoundFunction_STATE3[171]), .B(
        RoundFunction_T3_n591), .ZN(RoundFunction_TMP3_3[197]) );
  XNOR2_X1 RoundFunction_T3_U279 ( .A(RoundFunction_STATE3[170]), .B(
        RoundFunction_T3_n590), .ZN(RoundFunction_TMP3_3[196]) );
  XNOR2_X1 RoundFunction_T3_U278 ( .A(RoundFunction_STATE3[16]), .B(
        RoundFunction_T3_n596), .ZN(RoundFunction_TMP3_3[166]) );
  XNOR2_X1 RoundFunction_T3_U277 ( .A(RoundFunction_STATE3[169]), .B(
        RoundFunction_T3_n600), .ZN(RoundFunction_TMP3_3[195]) );
  XNOR2_X1 RoundFunction_T3_U276 ( .A(RoundFunction_STATE3[168]), .B(
        RoundFunction_T3_n589), .ZN(RoundFunction_TMP3_3[194]) );
  XNOR2_X1 RoundFunction_T3_U275 ( .A(RoundFunction_STATE3[167]), .B(
        RoundFunction_T3_n588), .ZN(RoundFunction_TMP3_3[113]) );
  XNOR2_X1 RoundFunction_T3_U274 ( .A(RoundFunction_STATE3[166]), .B(
        RoundFunction_T3_n587), .ZN(RoundFunction_TMP3_3[112]) );
  XNOR2_X1 RoundFunction_T3_U273 ( .A(RoundFunction_STATE3[165]), .B(
        RoundFunction_T3_n586), .ZN(RoundFunction_TMP3_3[119]) );
  XNOR2_X1 RoundFunction_T3_U272 ( .A(RoundFunction_STATE3[164]), .B(
        RoundFunction_T3_n585), .ZN(RoundFunction_TMP3_3[118]) );
  XNOR2_X1 RoundFunction_T3_U271 ( .A(RoundFunction_STATE3[163]), .B(
        RoundFunction_T3_n584), .ZN(RoundFunction_TMP3_3[117]) );
  XNOR2_X1 RoundFunction_T3_U270 ( .A(RoundFunction_STATE3[162]), .B(
        RoundFunction_T3_n583), .ZN(RoundFunction_TMP3_3[116]) );
  XNOR2_X1 RoundFunction_T3_U269 ( .A(RoundFunction_STATE3[161]), .B(
        RoundFunction_T3_n582), .ZN(RoundFunction_TMP3_3[115]) );
  XNOR2_X1 RoundFunction_T3_U268 ( .A(RoundFunction_STATE3[160]), .B(
        RoundFunction_T3_n581), .ZN(RoundFunction_TMP3_3[114]) );
  XNOR2_X1 RoundFunction_T3_U267 ( .A(RoundFunction_STATE3[15]), .B(
        RoundFunction_T3_n595), .ZN(RoundFunction_TMP3_3[80]) );
  XNOR2_X1 RoundFunction_T3_U266 ( .A(RoundFunction_STATE3[159]), .B(
        RoundFunction_T3_n580), .ZN(RoundFunction_TMP3_3[111]) );
  XNOR2_X1 RoundFunction_T3_U265 ( .A(RoundFunction_STATE3[158]), .B(
        RoundFunction_T3_n579), .ZN(RoundFunction_TMP3_3[110]) );
  XNOR2_X1 RoundFunction_T3_U264 ( .A(RoundFunction_STATE3[157]), .B(
        RoundFunction_T3_n578), .ZN(RoundFunction_TMP3_3[109]) );
  XNOR2_X1 RoundFunction_T3_U263 ( .A(RoundFunction_STATE3[156]), .B(
        RoundFunction_T3_n577), .ZN(RoundFunction_TMP3_3[108]) );
  XNOR2_X1 RoundFunction_T3_U262 ( .A(RoundFunction_STATE3[155]), .B(
        RoundFunction_T3_n576), .ZN(RoundFunction_TMP3_3[107]) );
  XNOR2_X1 RoundFunction_T3_U261 ( .A(RoundFunction_STATE3[154]), .B(
        RoundFunction_T3_n575), .ZN(RoundFunction_TMP3_3[106]) );
  XNOR2_X1 RoundFunction_T3_U260 ( .A(RoundFunction_STATE3[153]), .B(
        RoundFunction_T3_n574), .ZN(RoundFunction_TMP3_3[105]) );
  XNOR2_X1 RoundFunction_T3_U259 ( .A(RoundFunction_STATE3[152]), .B(
        RoundFunction_T3_n573), .ZN(RoundFunction_TMP3_3[104]) );
  XNOR2_X1 RoundFunction_T3_U258 ( .A(RoundFunction_STATE3[151]), .B(
        RoundFunction_T3_n572), .ZN(RoundFunction_TMP3_3[28]) );
  XNOR2_X1 RoundFunction_T3_U257 ( .A(RoundFunction_STATE3[150]), .B(
        RoundFunction_T3_n571), .ZN(RoundFunction_TMP3_3[27]) );
  XNOR2_X1 RoundFunction_T3_U256 ( .A(RoundFunction_STATE3[14]), .B(
        RoundFunction_T3_n594), .ZN(RoundFunction_TMP3_3[87]) );
  XNOR2_X1 RoundFunction_T3_U255 ( .A(RoundFunction_STATE3[149]), .B(
        RoundFunction_T3_n570), .ZN(RoundFunction_TMP3_3[26]) );
  XNOR2_X1 RoundFunction_T3_U254 ( .A(RoundFunction_STATE3[148]), .B(
        RoundFunction_T3_n569), .ZN(RoundFunction_TMP3_3[25]) );
  XNOR2_X1 RoundFunction_T3_U253 ( .A(RoundFunction_STATE3[147]), .B(
        RoundFunction_T3_n568), .ZN(RoundFunction_TMP3_3[24]) );
  XNOR2_X1 RoundFunction_T3_U252 ( .A(RoundFunction_STATE3[146]), .B(
        RoundFunction_T3_n567), .ZN(RoundFunction_TMP3_3[31]) );
  XNOR2_X1 RoundFunction_T3_U251 ( .A(RoundFunction_STATE3[145]), .B(
        RoundFunction_T3_n566), .ZN(RoundFunction_TMP3_3[30]) );
  XNOR2_X1 RoundFunction_T3_U250 ( .A(RoundFunction_STATE3[144]), .B(
        RoundFunction_T3_n565), .ZN(RoundFunction_TMP3_3[29]) );
  XNOR2_X1 RoundFunction_T3_U249 ( .A(RoundFunction_STATE3[143]), .B(
        RoundFunction_T3_n564), .ZN(RoundFunction_TMP3_3[150]) );
  XNOR2_X1 RoundFunction_T3_U248 ( .A(RoundFunction_STATE3[142]), .B(
        RoundFunction_T3_n563), .ZN(RoundFunction_TMP3_3[149]) );
  XNOR2_X1 RoundFunction_T3_U247 ( .A(RoundFunction_STATE3[141]), .B(
        RoundFunction_T3_n562), .ZN(RoundFunction_TMP3_3[148]) );
  XNOR2_X1 RoundFunction_T3_U246 ( .A(RoundFunction_STATE3[140]), .B(
        RoundFunction_T3_n561), .ZN(RoundFunction_TMP3_3[147]) );
  XNOR2_X1 RoundFunction_T3_U245 ( .A(RoundFunction_STATE3[13]), .B(
        RoundFunction_T3_n593), .ZN(RoundFunction_TMP3_3[86]) );
  XNOR2_X1 RoundFunction_T3_U244 ( .A(RoundFunction_STATE3[139]), .B(
        RoundFunction_T3_n599), .ZN(RoundFunction_TMP3_3[146]) );
  XNOR2_X1 RoundFunction_T3_U243 ( .A(RoundFunction_T3_n560), .B(
        RoundFunction_T3_n559), .ZN(RoundFunction_T3_n599) );
  XNOR2_X1 RoundFunction_T3_U242 ( .A(RoundFunction_STATE3[138]), .B(
        RoundFunction_T3_n598), .ZN(RoundFunction_TMP3_3[145]) );
  XNOR2_X1 RoundFunction_T3_U241 ( .A(RoundFunction_T3_n558), .B(
        RoundFunction_T3_n557), .ZN(RoundFunction_T3_n598) );
  XNOR2_X1 RoundFunction_T3_U240 ( .A(RoundFunction_STATE3[137]), .B(
        RoundFunction_T3_n597), .ZN(RoundFunction_TMP3_3[144]) );
  XNOR2_X1 RoundFunction_T3_U239 ( .A(RoundFunction_T3_n556), .B(
        RoundFunction_T3_n555), .ZN(RoundFunction_T3_n597) );
  XNOR2_X1 RoundFunction_T3_U238 ( .A(RoundFunction_STATE3[136]), .B(
        RoundFunction_T3_n596), .ZN(RoundFunction_TMP3_3[151]) );
  XNOR2_X1 RoundFunction_T3_U237 ( .A(RoundFunction_T3_n554), .B(
        RoundFunction_T3_n553), .ZN(RoundFunction_T3_n596) );
  XNOR2_X1 RoundFunction_T3_U236 ( .A(RoundFunction_STATE3[135]), .B(
        RoundFunction_T3_n595), .ZN(RoundFunction_TMP3_3[68]) );
  XNOR2_X1 RoundFunction_T3_U235 ( .A(RoundFunction_T3_n552), .B(
        RoundFunction_T3_n551), .ZN(RoundFunction_T3_n595) );
  XNOR2_X1 RoundFunction_T3_U234 ( .A(RoundFunction_STATE3[134]), .B(
        RoundFunction_T3_n594), .ZN(RoundFunction_TMP3_3[67]) );
  XNOR2_X1 RoundFunction_T3_U233 ( .A(RoundFunction_T3_n550), .B(
        RoundFunction_T3_n549), .ZN(RoundFunction_T3_n594) );
  XNOR2_X1 RoundFunction_T3_U232 ( .A(RoundFunction_STATE3[133]), .B(
        RoundFunction_T3_n593), .ZN(RoundFunction_TMP3_3[66]) );
  XNOR2_X1 RoundFunction_T3_U231 ( .A(RoundFunction_T3_n548), .B(
        RoundFunction_T3_n547), .ZN(RoundFunction_T3_n593) );
  XNOR2_X1 RoundFunction_T3_U230 ( .A(RoundFunction_STATE3[132]), .B(
        RoundFunction_T3_n592), .ZN(RoundFunction_TMP3_3[65]) );
  XNOR2_X1 RoundFunction_T3_U229 ( .A(RoundFunction_STATE3[131]), .B(
        RoundFunction_T3_n591), .ZN(RoundFunction_TMP3_3[64]) );
  XNOR2_X1 RoundFunction_T3_U228 ( .A(RoundFunction_STATE3[130]), .B(
        RoundFunction_T3_n590), .ZN(RoundFunction_TMP3_3[71]) );
  XNOR2_X1 RoundFunction_T3_U227 ( .A(RoundFunction_STATE3[12]), .B(
        RoundFunction_T3_n592), .ZN(RoundFunction_TMP3_3[85]) );
  XNOR2_X1 RoundFunction_T3_U226 ( .A(RoundFunction_T3_n546), .B(
        RoundFunction_T3_n545), .ZN(RoundFunction_T3_n592) );
  XNOR2_X1 RoundFunction_T3_U225 ( .A(RoundFunction_STATE3[129]), .B(
        RoundFunction_T3_n600), .ZN(RoundFunction_TMP3_3[70]) );
  XNOR2_X1 RoundFunction_T3_U224 ( .A(RoundFunction_T3_n544), .B(
        RoundFunction_T3_n543), .ZN(RoundFunction_T3_n600) );
  XNOR2_X1 RoundFunction_T3_U223 ( .A(RoundFunction_STATE3[128]), .B(
        RoundFunction_T3_n589), .ZN(RoundFunction_TMP3_3[69]) );
  XNOR2_X1 RoundFunction_T3_U222 ( .A(RoundFunction_T3_n542), .B(
        RoundFunction_T3_n541), .ZN(RoundFunction_T3_n589) );
  XNOR2_X1 RoundFunction_T3_U221 ( .A(RoundFunction_STATE3[127]), .B(
        RoundFunction_T3_n588), .ZN(RoundFunction_TMP3_3[184]) );
  XNOR2_X1 RoundFunction_T3_U220 ( .A(RoundFunction_T3_n540), .B(
        RoundFunction_T3_n539), .ZN(RoundFunction_T3_n588) );
  XNOR2_X1 RoundFunction_T3_U219 ( .A(RoundFunction_STATE3[126]), .B(
        RoundFunction_T3_n587), .ZN(RoundFunction_TMP3_3[191]) );
  XNOR2_X1 RoundFunction_T3_U218 ( .A(RoundFunction_T3_n538), .B(
        RoundFunction_T3_n537), .ZN(RoundFunction_T3_n587) );
  XNOR2_X1 RoundFunction_T3_U217 ( .A(RoundFunction_STATE3[125]), .B(
        RoundFunction_T3_n586), .ZN(RoundFunction_TMP3_3[190]) );
  XNOR2_X1 RoundFunction_T3_U216 ( .A(RoundFunction_T3_n536), .B(
        RoundFunction_T3_n535), .ZN(RoundFunction_T3_n586) );
  XNOR2_X1 RoundFunction_T3_U215 ( .A(RoundFunction_STATE3[124]), .B(
        RoundFunction_T3_n585), .ZN(RoundFunction_TMP3_3[189]) );
  XNOR2_X1 RoundFunction_T3_U214 ( .A(RoundFunction_T3_n534), .B(
        RoundFunction_T3_n559), .ZN(RoundFunction_T3_n585) );
  XOR2_X1 RoundFunction_T3_U213 ( .A(RoundFunction_STATE3[11]), .B(
        RoundFunction_T3_n533), .Z(RoundFunction_T3_n559) );
  XNOR2_X1 RoundFunction_T3_U212 ( .A(RoundFunction_T3_n532), .B(
        RoundFunction_T3_n531), .ZN(RoundFunction_T3_n533) );
  XNOR2_X1 RoundFunction_T3_U211 ( .A(RoundFunction_STATE3[51]), .B(
        RoundFunction_STATE3[91]), .ZN(RoundFunction_T3_n531) );
  XOR2_X1 RoundFunction_T3_U210 ( .A(RoundFunction_STATE3[131]), .B(
        RoundFunction_STATE3[171]), .Z(RoundFunction_T3_n532) );
  XNOR2_X1 RoundFunction_T3_U209 ( .A(RoundFunction_STATE3[123]), .B(
        RoundFunction_T3_n584), .ZN(RoundFunction_TMP3_3[188]) );
  XNOR2_X1 RoundFunction_T3_U208 ( .A(RoundFunction_T3_n530), .B(
        RoundFunction_T3_n557), .ZN(RoundFunction_T3_n584) );
  XOR2_X1 RoundFunction_T3_U207 ( .A(RoundFunction_STATE3[10]), .B(
        RoundFunction_T3_n529), .Z(RoundFunction_T3_n557) );
  XNOR2_X1 RoundFunction_T3_U206 ( .A(RoundFunction_T3_n528), .B(
        RoundFunction_T3_n527), .ZN(RoundFunction_T3_n529) );
  XNOR2_X1 RoundFunction_T3_U205 ( .A(RoundFunction_STATE3[50]), .B(
        RoundFunction_STATE3[90]), .ZN(RoundFunction_T3_n527) );
  XOR2_X1 RoundFunction_T3_U204 ( .A(RoundFunction_STATE3[130]), .B(
        RoundFunction_STATE3[170]), .Z(RoundFunction_T3_n528) );
  XNOR2_X1 RoundFunction_T3_U203 ( .A(RoundFunction_STATE3[122]), .B(
        RoundFunction_T3_n583), .ZN(RoundFunction_TMP3_3[187]) );
  XNOR2_X1 RoundFunction_T3_U202 ( .A(RoundFunction_T3_n526), .B(
        RoundFunction_T3_n555), .ZN(RoundFunction_T3_n583) );
  XOR2_X1 RoundFunction_T3_U201 ( .A(RoundFunction_STATE3[89]), .B(
        RoundFunction_T3_n525), .Z(RoundFunction_T3_n555) );
  XNOR2_X1 RoundFunction_T3_U200 ( .A(RoundFunction_T3_n524), .B(
        RoundFunction_T3_n523), .ZN(RoundFunction_T3_n525) );
  XNOR2_X1 RoundFunction_T3_U199 ( .A(RoundFunction_STATE3[129]), .B(
        RoundFunction_STATE3[49]), .ZN(RoundFunction_T3_n523) );
  XOR2_X1 RoundFunction_T3_U198 ( .A(RoundFunction_STATE3[169]), .B(
        RoundFunction_STATE3[9]), .Z(RoundFunction_T3_n524) );
  XNOR2_X1 RoundFunction_T3_U197 ( .A(RoundFunction_STATE3[121]), .B(
        RoundFunction_T3_n582), .ZN(RoundFunction_TMP3_3[186]) );
  XNOR2_X1 RoundFunction_T3_U196 ( .A(RoundFunction_T3_n522), .B(
        RoundFunction_T3_n553), .ZN(RoundFunction_T3_n582) );
  XOR2_X1 RoundFunction_T3_U195 ( .A(RoundFunction_STATE3[128]), .B(
        RoundFunction_T3_n521), .Z(RoundFunction_T3_n553) );
  XNOR2_X1 RoundFunction_T3_U194 ( .A(RoundFunction_T3_n520), .B(
        RoundFunction_T3_n519), .ZN(RoundFunction_T3_n521) );
  XNOR2_X1 RoundFunction_T3_U193 ( .A(RoundFunction_STATE3[48]), .B(
        RoundFunction_STATE3[8]), .ZN(RoundFunction_T3_n519) );
  XOR2_X1 RoundFunction_T3_U192 ( .A(RoundFunction_STATE3[88]), .B(
        RoundFunction_STATE3[168]), .Z(RoundFunction_T3_n520) );
  XNOR2_X1 RoundFunction_T3_U191 ( .A(RoundFunction_STATE3[120]), .B(
        RoundFunction_T3_n581), .ZN(RoundFunction_TMP3_3[185]) );
  XNOR2_X1 RoundFunction_T3_U190 ( .A(RoundFunction_STATE3[11]), .B(
        RoundFunction_T3_n591), .ZN(RoundFunction_TMP3_3[84]) );
  XNOR2_X1 RoundFunction_T3_U189 ( .A(RoundFunction_T3_n518), .B(
        RoundFunction_T3_n517), .ZN(RoundFunction_T3_n591) );
  XNOR2_X1 RoundFunction_T3_U188 ( .A(RoundFunction_STATE3[119]), .B(
        RoundFunction_T3_n580), .ZN(RoundFunction_TMP3_3[182]) );
  XNOR2_X1 RoundFunction_T3_U187 ( .A(RoundFunction_T3_n554), .B(
        RoundFunction_T3_n549), .ZN(RoundFunction_T3_n580) );
  XOR2_X1 RoundFunction_T3_U186 ( .A(RoundFunction_STATE3[126]), .B(
        RoundFunction_T3_n516), .Z(RoundFunction_T3_n549) );
  XNOR2_X1 RoundFunction_T3_U185 ( .A(RoundFunction_T3_n515), .B(
        RoundFunction_T3_n514), .ZN(RoundFunction_T3_n516) );
  XNOR2_X1 RoundFunction_T3_U184 ( .A(RoundFunction_STATE3[46]), .B(
        RoundFunction_STATE3[86]), .ZN(RoundFunction_T3_n514) );
  XOR2_X1 RoundFunction_T3_U183 ( .A(RoundFunction_STATE3[6]), .B(
        RoundFunction_STATE3[166]), .Z(RoundFunction_T3_n515) );
  XOR2_X1 RoundFunction_T3_U182 ( .A(RoundFunction_STATE3[111]), .B(
        RoundFunction_T3_n513), .Z(RoundFunction_T3_n554) );
  XNOR2_X1 RoundFunction_T3_U181 ( .A(RoundFunction_T3_n512), .B(
        RoundFunction_T3_n511), .ZN(RoundFunction_T3_n513) );
  XNOR2_X1 RoundFunction_T3_U180 ( .A(RoundFunction_STATE3[31]), .B(
        RoundFunction_STATE3[71]), .ZN(RoundFunction_T3_n511) );
  XOR2_X1 RoundFunction_T3_U179 ( .A(RoundFunction_STATE3[151]), .B(
        RoundFunction_STATE3[191]), .Z(RoundFunction_T3_n512) );
  XNOR2_X1 RoundFunction_T3_U178 ( .A(RoundFunction_STATE3[118]), .B(
        RoundFunction_T3_n579), .ZN(RoundFunction_TMP3_3[181]) );
  XNOR2_X1 RoundFunction_T3_U177 ( .A(RoundFunction_T3_n510), .B(
        RoundFunction_T3_n547), .ZN(RoundFunction_T3_n579) );
  XOR2_X1 RoundFunction_T3_U176 ( .A(RoundFunction_STATE3[125]), .B(
        RoundFunction_T3_n509), .Z(RoundFunction_T3_n547) );
  XNOR2_X1 RoundFunction_T3_U175 ( .A(RoundFunction_T3_n508), .B(
        RoundFunction_T3_n507), .ZN(RoundFunction_T3_n509) );
  XNOR2_X1 RoundFunction_T3_U174 ( .A(RoundFunction_STATE3[45]), .B(
        RoundFunction_STATE3[85]), .ZN(RoundFunction_T3_n507) );
  XOR2_X1 RoundFunction_T3_U173 ( .A(RoundFunction_STATE3[5]), .B(
        RoundFunction_STATE3[165]), .Z(RoundFunction_T3_n508) );
  XNOR2_X1 RoundFunction_T3_U172 ( .A(RoundFunction_STATE3[117]), .B(
        RoundFunction_T3_n578), .ZN(RoundFunction_TMP3_3[180]) );
  XNOR2_X1 RoundFunction_T3_U171 ( .A(RoundFunction_T3_n506), .B(
        RoundFunction_T3_n545), .ZN(RoundFunction_T3_n578) );
  XOR2_X1 RoundFunction_T3_U170 ( .A(RoundFunction_STATE3[124]), .B(
        RoundFunction_T3_n505), .Z(RoundFunction_T3_n545) );
  XNOR2_X1 RoundFunction_T3_U169 ( .A(RoundFunction_T3_n504), .B(
        RoundFunction_T3_n503), .ZN(RoundFunction_T3_n505) );
  XNOR2_X1 RoundFunction_T3_U168 ( .A(RoundFunction_STATE3[44]), .B(
        RoundFunction_STATE3[84]), .ZN(RoundFunction_T3_n503) );
  XOR2_X1 RoundFunction_T3_U167 ( .A(RoundFunction_STATE3[4]), .B(
        RoundFunction_STATE3[164]), .Z(RoundFunction_T3_n504) );
  XNOR2_X1 RoundFunction_T3_U166 ( .A(RoundFunction_STATE3[116]), .B(
        RoundFunction_T3_n577), .ZN(RoundFunction_TMP3_3[179]) );
  XNOR2_X1 RoundFunction_T3_U165 ( .A(RoundFunction_T3_n502), .B(
        RoundFunction_T3_n517), .ZN(RoundFunction_T3_n577) );
  XOR2_X1 RoundFunction_T3_U164 ( .A(RoundFunction_STATE3[123]), .B(
        RoundFunction_T3_n501), .Z(RoundFunction_T3_n517) );
  XNOR2_X1 RoundFunction_T3_U163 ( .A(RoundFunction_T3_n500), .B(
        RoundFunction_T3_n499), .ZN(RoundFunction_T3_n501) );
  XNOR2_X1 RoundFunction_T3_U162 ( .A(RoundFunction_STATE3[3]), .B(
        RoundFunction_STATE3[83]), .ZN(RoundFunction_T3_n499) );
  XOR2_X1 RoundFunction_T3_U161 ( .A(RoundFunction_STATE3[43]), .B(
        RoundFunction_STATE3[163]), .Z(RoundFunction_T3_n500) );
  XNOR2_X1 RoundFunction_T3_U160 ( .A(RoundFunction_STATE3[115]), .B(
        RoundFunction_T3_n576), .ZN(RoundFunction_TMP3_3[178]) );
  XNOR2_X1 RoundFunction_T3_U159 ( .A(RoundFunction_T3_n498), .B(
        RoundFunction_T3_n497), .ZN(RoundFunction_T3_n576) );
  XNOR2_X1 RoundFunction_T3_U158 ( .A(RoundFunction_STATE3[114]), .B(
        RoundFunction_T3_n575), .ZN(RoundFunction_TMP3_3[177]) );
  XNOR2_X1 RoundFunction_T3_U157 ( .A(RoundFunction_T3_n543), .B(
        RoundFunction_T3_n560), .ZN(RoundFunction_T3_n575) );
  XOR2_X1 RoundFunction_T3_U156 ( .A(RoundFunction_STATE3[106]), .B(
        RoundFunction_T3_n496), .Z(RoundFunction_T3_n560) );
  XNOR2_X1 RoundFunction_T3_U155 ( .A(RoundFunction_T3_n495), .B(
        RoundFunction_T3_n494), .ZN(RoundFunction_T3_n496) );
  XNOR2_X1 RoundFunction_T3_U154 ( .A(RoundFunction_STATE3[26]), .B(
        RoundFunction_STATE3[66]), .ZN(RoundFunction_T3_n494) );
  XOR2_X1 RoundFunction_T3_U153 ( .A(RoundFunction_STATE3[146]), .B(
        RoundFunction_STATE3[186]), .Z(RoundFunction_T3_n495) );
  XOR2_X1 RoundFunction_T3_U152 ( .A(RoundFunction_STATE3[121]), .B(
        RoundFunction_T3_n493), .Z(RoundFunction_T3_n543) );
  XNOR2_X1 RoundFunction_T3_U151 ( .A(RoundFunction_T3_n492), .B(
        RoundFunction_T3_n491), .ZN(RoundFunction_T3_n493) );
  XNOR2_X1 RoundFunction_T3_U150 ( .A(RoundFunction_STATE3[1]), .B(
        RoundFunction_STATE3[81]), .ZN(RoundFunction_T3_n491) );
  XOR2_X1 RoundFunction_T3_U149 ( .A(RoundFunction_STATE3[41]), .B(
        RoundFunction_STATE3[161]), .Z(RoundFunction_T3_n492) );
  XNOR2_X1 RoundFunction_T3_U148 ( .A(RoundFunction_STATE3[113]), .B(
        RoundFunction_T3_n574), .ZN(RoundFunction_TMP3_3[176]) );
  XNOR2_X1 RoundFunction_T3_U147 ( .A(RoundFunction_T3_n558), .B(
        RoundFunction_T3_n541), .ZN(RoundFunction_T3_n574) );
  XOR2_X1 RoundFunction_T3_U146 ( .A(RoundFunction_STATE3[0]), .B(
        RoundFunction_T3_n490), .Z(RoundFunction_T3_n541) );
  XNOR2_X1 RoundFunction_T3_U145 ( .A(RoundFunction_T3_n489), .B(
        RoundFunction_T3_n488), .ZN(RoundFunction_T3_n490) );
  XNOR2_X1 RoundFunction_T3_U144 ( .A(RoundFunction_STATE3[40]), .B(
        RoundFunction_STATE3[80]), .ZN(RoundFunction_T3_n488) );
  XOR2_X1 RoundFunction_T3_U143 ( .A(RoundFunction_STATE3[120]), .B(
        RoundFunction_STATE3[160]), .Z(RoundFunction_T3_n489) );
  XOR2_X1 RoundFunction_T3_U142 ( .A(RoundFunction_STATE3[105]), .B(
        RoundFunction_T3_n487), .Z(RoundFunction_T3_n558) );
  XNOR2_X1 RoundFunction_T3_U141 ( .A(RoundFunction_T3_n486), .B(
        RoundFunction_T3_n485), .ZN(RoundFunction_T3_n487) );
  XNOR2_X1 RoundFunction_T3_U140 ( .A(RoundFunction_STATE3[25]), .B(
        RoundFunction_STATE3[65]), .ZN(RoundFunction_T3_n485) );
  XOR2_X1 RoundFunction_T3_U139 ( .A(RoundFunction_STATE3[145]), .B(
        RoundFunction_STATE3[185]), .Z(RoundFunction_T3_n486) );
  XNOR2_X1 RoundFunction_T3_U138 ( .A(RoundFunction_STATE3[112]), .B(
        RoundFunction_T3_n573), .ZN(RoundFunction_TMP3_3[183]) );
  XNOR2_X1 RoundFunction_T3_U137 ( .A(RoundFunction_T3_n556), .B(
        RoundFunction_T3_n551), .ZN(RoundFunction_T3_n573) );
  XOR2_X1 RoundFunction_T3_U136 ( .A(RoundFunction_STATE3[127]), .B(
        RoundFunction_T3_n484), .Z(RoundFunction_T3_n551) );
  XNOR2_X1 RoundFunction_T3_U135 ( .A(RoundFunction_T3_n483), .B(
        RoundFunction_T3_n482), .ZN(RoundFunction_T3_n484) );
  XNOR2_X1 RoundFunction_T3_U134 ( .A(RoundFunction_STATE3[47]), .B(
        RoundFunction_STATE3[87]), .ZN(RoundFunction_T3_n482) );
  XOR2_X1 RoundFunction_T3_U133 ( .A(RoundFunction_STATE3[7]), .B(
        RoundFunction_STATE3[167]), .Z(RoundFunction_T3_n483) );
  XOR2_X1 RoundFunction_T3_U132 ( .A(RoundFunction_STATE3[104]), .B(
        RoundFunction_T3_n481), .Z(RoundFunction_T3_n556) );
  XNOR2_X1 RoundFunction_T3_U131 ( .A(RoundFunction_T3_n480), .B(
        RoundFunction_T3_n479), .ZN(RoundFunction_T3_n481) );
  XNOR2_X1 RoundFunction_T3_U130 ( .A(RoundFunction_STATE3[24]), .B(
        RoundFunction_STATE3[64]), .ZN(RoundFunction_T3_n479) );
  XOR2_X1 RoundFunction_T3_U129 ( .A(RoundFunction_STATE3[144]), .B(
        RoundFunction_STATE3[184]), .Z(RoundFunction_T3_n480) );
  XNOR2_X1 RoundFunction_T3_U128 ( .A(RoundFunction_STATE3[111]), .B(
        RoundFunction_T3_n572), .ZN(RoundFunction_TMP3_3[96]) );
  XNOR2_X1 RoundFunction_T3_U127 ( .A(RoundFunction_T3_n542), .B(
        RoundFunction_T3_n537), .ZN(RoundFunction_T3_n572) );
  XOR2_X1 RoundFunction_T3_U126 ( .A(RoundFunction_STATE3[118]), .B(
        RoundFunction_T3_n478), .Z(RoundFunction_T3_n537) );
  XNOR2_X1 RoundFunction_T3_U125 ( .A(RoundFunction_T3_n477), .B(
        RoundFunction_T3_n476), .ZN(RoundFunction_T3_n478) );
  XNOR2_X1 RoundFunction_T3_U124 ( .A(RoundFunction_STATE3[198]), .B(
        RoundFunction_STATE3[78]), .ZN(RoundFunction_T3_n476) );
  XOR2_X1 RoundFunction_T3_U123 ( .A(RoundFunction_STATE3[38]), .B(
        RoundFunction_STATE3[158]), .Z(RoundFunction_T3_n477) );
  XOR2_X1 RoundFunction_T3_U122 ( .A(RoundFunction_STATE3[103]), .B(
        RoundFunction_T3_n475), .Z(RoundFunction_T3_n542) );
  XNOR2_X1 RoundFunction_T3_U121 ( .A(RoundFunction_T3_n474), .B(
        RoundFunction_T3_n473), .ZN(RoundFunction_T3_n475) );
  XNOR2_X1 RoundFunction_T3_U120 ( .A(RoundFunction_STATE3[23]), .B(
        RoundFunction_STATE3[63]), .ZN(RoundFunction_T3_n473) );
  XOR2_X1 RoundFunction_T3_U119 ( .A(RoundFunction_STATE3[143]), .B(
        RoundFunction_STATE3[183]), .Z(RoundFunction_T3_n474) );
  XNOR2_X1 RoundFunction_T3_U118 ( .A(RoundFunction_STATE3[110]), .B(
        RoundFunction_T3_n571), .ZN(RoundFunction_TMP3_3[103]) );
  XNOR2_X1 RoundFunction_T3_U117 ( .A(RoundFunction_T3_n552), .B(
        RoundFunction_T3_n535), .ZN(RoundFunction_T3_n571) );
  XOR2_X1 RoundFunction_T3_U116 ( .A(RoundFunction_STATE3[117]), .B(
        RoundFunction_T3_n472), .Z(RoundFunction_T3_n535) );
  XNOR2_X1 RoundFunction_T3_U115 ( .A(RoundFunction_T3_n471), .B(
        RoundFunction_T3_n470), .ZN(RoundFunction_T3_n472) );
  XNOR2_X1 RoundFunction_T3_U114 ( .A(RoundFunction_STATE3[197]), .B(
        RoundFunction_STATE3[77]), .ZN(RoundFunction_T3_n470) );
  XOR2_X1 RoundFunction_T3_U113 ( .A(RoundFunction_STATE3[37]), .B(
        RoundFunction_STATE3[157]), .Z(RoundFunction_T3_n471) );
  XOR2_X1 RoundFunction_T3_U112 ( .A(RoundFunction_STATE3[102]), .B(
        RoundFunction_T3_n469), .Z(RoundFunction_T3_n552) );
  XNOR2_X1 RoundFunction_T3_U111 ( .A(RoundFunction_T3_n468), .B(
        RoundFunction_T3_n467), .ZN(RoundFunction_T3_n469) );
  XNOR2_X1 RoundFunction_T3_U110 ( .A(RoundFunction_STATE3[22]), .B(
        RoundFunction_STATE3[62]), .ZN(RoundFunction_T3_n467) );
  XOR2_X1 RoundFunction_T3_U109 ( .A(RoundFunction_STATE3[142]), .B(
        RoundFunction_STATE3[182]), .Z(RoundFunction_T3_n468) );
  XNOR2_X1 RoundFunction_T3_U108 ( .A(RoundFunction_STATE3[10]), .B(
        RoundFunction_T3_n590), .ZN(RoundFunction_TMP3_3[83]) );
  XNOR2_X1 RoundFunction_T3_U107 ( .A(RoundFunction_T3_n466), .B(
        RoundFunction_T3_n497), .ZN(RoundFunction_T3_n590) );
  XOR2_X1 RoundFunction_T3_U106 ( .A(RoundFunction_STATE3[122]), .B(
        RoundFunction_T3_n465), .Z(RoundFunction_T3_n497) );
  XNOR2_X1 RoundFunction_T3_U105 ( .A(RoundFunction_T3_n464), .B(
        RoundFunction_T3_n463), .ZN(RoundFunction_T3_n465) );
  XNOR2_X1 RoundFunction_T3_U104 ( .A(RoundFunction_STATE3[2]), .B(
        RoundFunction_STATE3[82]), .ZN(RoundFunction_T3_n463) );
  XOR2_X1 RoundFunction_T3_U103 ( .A(RoundFunction_STATE3[42]), .B(
        RoundFunction_STATE3[162]), .Z(RoundFunction_T3_n464) );
  XNOR2_X1 RoundFunction_T3_U102 ( .A(RoundFunction_STATE3[109]), .B(
        RoundFunction_T3_n570), .ZN(RoundFunction_TMP3_3[102]) );
  XNOR2_X1 RoundFunction_T3_U101 ( .A(RoundFunction_T3_n550), .B(
        RoundFunction_T3_n534), .ZN(RoundFunction_T3_n570) );
  XOR2_X1 RoundFunction_T3_U100 ( .A(RoundFunction_STATE3[116]), .B(
        RoundFunction_T3_n462), .Z(RoundFunction_T3_n534) );
  XNOR2_X1 RoundFunction_T3_U99 ( .A(RoundFunction_T3_n461), .B(
        RoundFunction_T3_n460), .ZN(RoundFunction_T3_n462) );
  XNOR2_X1 RoundFunction_T3_U98 ( .A(RoundFunction_STATE3[196]), .B(
        RoundFunction_STATE3[76]), .ZN(RoundFunction_T3_n460) );
  XOR2_X1 RoundFunction_T3_U97 ( .A(RoundFunction_STATE3[36]), .B(
        RoundFunction_STATE3[156]), .Z(RoundFunction_T3_n461) );
  XOR2_X1 RoundFunction_T3_U96 ( .A(RoundFunction_STATE3[101]), .B(
        RoundFunction_T3_n459), .Z(RoundFunction_T3_n550) );
  XNOR2_X1 RoundFunction_T3_U95 ( .A(RoundFunction_T3_n458), .B(
        RoundFunction_T3_n457), .ZN(RoundFunction_T3_n459) );
  XNOR2_X1 RoundFunction_T3_U94 ( .A(RoundFunction_STATE3[21]), .B(
        RoundFunction_STATE3[61]), .ZN(RoundFunction_T3_n457) );
  XOR2_X1 RoundFunction_T3_U93 ( .A(RoundFunction_STATE3[141]), .B(
        RoundFunction_STATE3[181]), .Z(RoundFunction_T3_n458) );
  XNOR2_X1 RoundFunction_T3_U92 ( .A(RoundFunction_STATE3[108]), .B(
        RoundFunction_T3_n569), .ZN(RoundFunction_TMP3_3[101]) );
  XNOR2_X1 RoundFunction_T3_U91 ( .A(RoundFunction_T3_n548), .B(
        RoundFunction_T3_n530), .ZN(RoundFunction_T3_n569) );
  XOR2_X1 RoundFunction_T3_U90 ( .A(RoundFunction_STATE3[115]), .B(
        RoundFunction_T3_n456), .Z(RoundFunction_T3_n530) );
  XNOR2_X1 RoundFunction_T3_U89 ( .A(RoundFunction_T3_n455), .B(
        RoundFunction_T3_n454), .ZN(RoundFunction_T3_n456) );
  XNOR2_X1 RoundFunction_T3_U88 ( .A(RoundFunction_STATE3[195]), .B(
        RoundFunction_STATE3[75]), .ZN(RoundFunction_T3_n454) );
  XOR2_X1 RoundFunction_T3_U87 ( .A(RoundFunction_STATE3[35]), .B(
        RoundFunction_STATE3[155]), .Z(RoundFunction_T3_n455) );
  XOR2_X1 RoundFunction_T3_U86 ( .A(RoundFunction_STATE3[100]), .B(
        RoundFunction_T3_n453), .Z(RoundFunction_T3_n548) );
  XNOR2_X1 RoundFunction_T3_U85 ( .A(RoundFunction_T3_n452), .B(
        RoundFunction_T3_n451), .ZN(RoundFunction_T3_n453) );
  XNOR2_X1 RoundFunction_T3_U84 ( .A(RoundFunction_STATE3[20]), .B(
        RoundFunction_STATE3[60]), .ZN(RoundFunction_T3_n451) );
  XOR2_X1 RoundFunction_T3_U83 ( .A(RoundFunction_STATE3[140]), .B(
        RoundFunction_STATE3[180]), .Z(RoundFunction_T3_n452) );
  XNOR2_X1 RoundFunction_T3_U82 ( .A(RoundFunction_STATE3[107]), .B(
        RoundFunction_T3_n568), .ZN(RoundFunction_TMP3_3[100]) );
  XNOR2_X1 RoundFunction_T3_U81 ( .A(RoundFunction_T3_n546), .B(
        RoundFunction_T3_n526), .ZN(RoundFunction_T3_n568) );
  XOR2_X1 RoundFunction_T3_U80 ( .A(RoundFunction_STATE3[114]), .B(
        RoundFunction_T3_n450), .Z(RoundFunction_T3_n526) );
  XNOR2_X1 RoundFunction_T3_U79 ( .A(RoundFunction_T3_n449), .B(
        RoundFunction_T3_n448), .ZN(RoundFunction_T3_n450) );
  XNOR2_X1 RoundFunction_T3_U78 ( .A(RoundFunction_STATE3[194]), .B(
        RoundFunction_STATE3[74]), .ZN(RoundFunction_T3_n448) );
  XOR2_X1 RoundFunction_T3_U77 ( .A(RoundFunction_STATE3[34]), .B(
        RoundFunction_STATE3[154]), .Z(RoundFunction_T3_n449) );
  XOR2_X1 RoundFunction_T3_U76 ( .A(RoundFunction_STATE3[59]), .B(
        RoundFunction_T3_n447), .Z(RoundFunction_T3_n546) );
  XNOR2_X1 RoundFunction_T3_U75 ( .A(RoundFunction_T3_n446), .B(
        RoundFunction_T3_n445), .ZN(RoundFunction_T3_n447) );
  XNOR2_X1 RoundFunction_T3_U74 ( .A(RoundFunction_STATE3[139]), .B(
        RoundFunction_STATE3[19]), .ZN(RoundFunction_T3_n445) );
  XOR2_X1 RoundFunction_T3_U73 ( .A(RoundFunction_STATE3[179]), .B(
        RoundFunction_STATE3[99]), .Z(RoundFunction_T3_n446) );
  XNOR2_X1 RoundFunction_T3_U72 ( .A(RoundFunction_STATE3[106]), .B(
        RoundFunction_T3_n567), .ZN(RoundFunction_TMP3_3[99]) );
  XNOR2_X1 RoundFunction_T3_U71 ( .A(RoundFunction_T3_n518), .B(
        RoundFunction_T3_n522), .ZN(RoundFunction_T3_n567) );
  XOR2_X1 RoundFunction_T3_U70 ( .A(RoundFunction_STATE3[113]), .B(
        RoundFunction_T3_n444), .Z(RoundFunction_T3_n522) );
  XNOR2_X1 RoundFunction_T3_U69 ( .A(RoundFunction_T3_n443), .B(
        RoundFunction_T3_n442), .ZN(RoundFunction_T3_n444) );
  XNOR2_X1 RoundFunction_T3_U68 ( .A(RoundFunction_STATE3[193]), .B(
        RoundFunction_STATE3[73]), .ZN(RoundFunction_T3_n442) );
  XOR2_X1 RoundFunction_T3_U67 ( .A(RoundFunction_STATE3[33]), .B(
        RoundFunction_STATE3[153]), .Z(RoundFunction_T3_n443) );
  XOR2_X1 RoundFunction_T3_U66 ( .A(RoundFunction_STATE3[58]), .B(
        RoundFunction_T3_n441), .Z(RoundFunction_T3_n518) );
  XNOR2_X1 RoundFunction_T3_U65 ( .A(RoundFunction_T3_n440), .B(
        RoundFunction_T3_n439), .ZN(RoundFunction_T3_n441) );
  XNOR2_X1 RoundFunction_T3_U64 ( .A(RoundFunction_STATE3[138]), .B(
        RoundFunction_STATE3[18]), .ZN(RoundFunction_T3_n439) );
  XOR2_X1 RoundFunction_T3_U63 ( .A(RoundFunction_STATE3[178]), .B(
        RoundFunction_STATE3[98]), .Z(RoundFunction_T3_n440) );
  XNOR2_X1 RoundFunction_T3_U62 ( .A(RoundFunction_STATE3[105]), .B(
        RoundFunction_T3_n566), .ZN(RoundFunction_TMP3_3[98]) );
  XNOR2_X1 RoundFunction_T3_U61 ( .A(RoundFunction_T3_n438), .B(
        RoundFunction_T3_n466), .ZN(RoundFunction_T3_n566) );
  XOR2_X1 RoundFunction_T3_U60 ( .A(RoundFunction_STATE3[57]), .B(
        RoundFunction_T3_n437), .Z(RoundFunction_T3_n466) );
  XNOR2_X1 RoundFunction_T3_U59 ( .A(RoundFunction_T3_n436), .B(
        RoundFunction_T3_n435), .ZN(RoundFunction_T3_n437) );
  XNOR2_X1 RoundFunction_T3_U58 ( .A(RoundFunction_STATE3[137]), .B(
        RoundFunction_STATE3[17]), .ZN(RoundFunction_T3_n435) );
  XOR2_X1 RoundFunction_T3_U57 ( .A(RoundFunction_STATE3[177]), .B(
        RoundFunction_STATE3[97]), .Z(RoundFunction_T3_n436) );
  XNOR2_X1 RoundFunction_T3_U56 ( .A(RoundFunction_STATE3[104]), .B(
        RoundFunction_T3_n565), .ZN(RoundFunction_TMP3_3[97]) );
  XNOR2_X1 RoundFunction_T3_U55 ( .A(RoundFunction_T3_n544), .B(
        RoundFunction_T3_n539), .ZN(RoundFunction_T3_n565) );
  XOR2_X1 RoundFunction_T3_U54 ( .A(RoundFunction_STATE3[119]), .B(
        RoundFunction_T3_n434), .Z(RoundFunction_T3_n539) );
  XNOR2_X1 RoundFunction_T3_U53 ( .A(RoundFunction_T3_n433), .B(
        RoundFunction_T3_n432), .ZN(RoundFunction_T3_n434) );
  XNOR2_X1 RoundFunction_T3_U52 ( .A(RoundFunction_STATE3[199]), .B(
        RoundFunction_STATE3[79]), .ZN(RoundFunction_T3_n432) );
  XOR2_X1 RoundFunction_T3_U51 ( .A(RoundFunction_STATE3[39]), .B(
        RoundFunction_STATE3[159]), .Z(RoundFunction_T3_n433) );
  XOR2_X1 RoundFunction_T3_U50 ( .A(RoundFunction_STATE3[136]), .B(
        RoundFunction_T3_n431), .Z(RoundFunction_T3_n544) );
  XNOR2_X1 RoundFunction_T3_U49 ( .A(RoundFunction_T3_n430), .B(
        RoundFunction_T3_n429), .ZN(RoundFunction_T3_n431) );
  XNOR2_X1 RoundFunction_T3_U48 ( .A(RoundFunction_STATE3[176]), .B(
        RoundFunction_STATE3[96]), .ZN(RoundFunction_T3_n429) );
  XOR2_X1 RoundFunction_T3_U47 ( .A(RoundFunction_STATE3[56]), .B(
        RoundFunction_STATE3[16]), .Z(RoundFunction_T3_n430) );
  XNOR2_X1 RoundFunction_T3_U46 ( .A(RoundFunction_STATE3[103]), .B(
        RoundFunction_T3_n564), .ZN(RoundFunction_TMP3_3[18]) );
  XNOR2_X1 RoundFunction_T3_U45 ( .A(RoundFunction_T3_n428), .B(
        RoundFunction_T3_n510), .ZN(RoundFunction_T3_n564) );
  XOR2_X1 RoundFunction_T3_U44 ( .A(RoundFunction_STATE3[110]), .B(
        RoundFunction_T3_n427), .Z(RoundFunction_T3_n510) );
  XNOR2_X1 RoundFunction_T3_U43 ( .A(RoundFunction_T3_n426), .B(
        RoundFunction_T3_n425), .ZN(RoundFunction_T3_n427) );
  XNOR2_X1 RoundFunction_T3_U42 ( .A(RoundFunction_STATE3[190]), .B(
        RoundFunction_STATE3[70]), .ZN(RoundFunction_T3_n425) );
  XOR2_X1 RoundFunction_T3_U41 ( .A(RoundFunction_STATE3[30]), .B(
        RoundFunction_STATE3[150]), .Z(RoundFunction_T3_n426) );
  XNOR2_X1 RoundFunction_T3_U40 ( .A(RoundFunction_STATE3[102]), .B(
        RoundFunction_T3_n563), .ZN(RoundFunction_TMP3_3[17]) );
  XNOR2_X1 RoundFunction_T3_U39 ( .A(RoundFunction_T3_n540), .B(
        RoundFunction_T3_n506), .ZN(RoundFunction_T3_n563) );
  XOR2_X1 RoundFunction_T3_U38 ( .A(RoundFunction_STATE3[109]), .B(
        RoundFunction_T3_n424), .Z(RoundFunction_T3_n506) );
  XNOR2_X1 RoundFunction_T3_U37 ( .A(RoundFunction_T3_n423), .B(
        RoundFunction_T3_n422), .ZN(RoundFunction_T3_n424) );
  XNOR2_X1 RoundFunction_T3_U36 ( .A(RoundFunction_STATE3[189]), .B(
        RoundFunction_STATE3[69]), .ZN(RoundFunction_T3_n422) );
  XOR2_X1 RoundFunction_T3_U35 ( .A(RoundFunction_STATE3[29]), .B(
        RoundFunction_STATE3[149]), .Z(RoundFunction_T3_n423) );
  XOR2_X1 RoundFunction_T3_U34 ( .A(RoundFunction_STATE3[54]), .B(
        RoundFunction_T3_n421), .Z(RoundFunction_T3_n540) );
  XNOR2_X1 RoundFunction_T3_U33 ( .A(RoundFunction_T3_n420), .B(
        RoundFunction_T3_n419), .ZN(RoundFunction_T3_n421) );
  XNOR2_X1 RoundFunction_T3_U32 ( .A(RoundFunction_STATE3[134]), .B(
        RoundFunction_STATE3[174]), .ZN(RoundFunction_T3_n419) );
  XOR2_X1 RoundFunction_T3_U31 ( .A(RoundFunction_STATE3[14]), .B(
        RoundFunction_STATE3[94]), .Z(RoundFunction_T3_n420) );
  XNOR2_X1 RoundFunction_T3_U30 ( .A(RoundFunction_STATE3[101]), .B(
        RoundFunction_T3_n562), .ZN(RoundFunction_TMP3_3[16]) );
  XNOR2_X1 RoundFunction_T3_U29 ( .A(RoundFunction_T3_n538), .B(
        RoundFunction_T3_n502), .ZN(RoundFunction_T3_n562) );
  XOR2_X1 RoundFunction_T3_U28 ( .A(RoundFunction_STATE3[108]), .B(
        RoundFunction_T3_n418), .Z(RoundFunction_T3_n502) );
  XNOR2_X1 RoundFunction_T3_U27 ( .A(RoundFunction_T3_n417), .B(
        RoundFunction_T3_n416), .ZN(RoundFunction_T3_n418) );
  XNOR2_X1 RoundFunction_T3_U26 ( .A(RoundFunction_STATE3[188]), .B(
        RoundFunction_STATE3[68]), .ZN(RoundFunction_T3_n416) );
  XOR2_X1 RoundFunction_T3_U25 ( .A(RoundFunction_STATE3[28]), .B(
        RoundFunction_STATE3[148]), .Z(RoundFunction_T3_n417) );
  XOR2_X1 RoundFunction_T3_U24 ( .A(RoundFunction_STATE3[53]), .B(
        RoundFunction_T3_n415), .Z(RoundFunction_T3_n538) );
  XNOR2_X1 RoundFunction_T3_U23 ( .A(RoundFunction_T3_n414), .B(
        RoundFunction_T3_n413), .ZN(RoundFunction_T3_n415) );
  XNOR2_X1 RoundFunction_T3_U22 ( .A(RoundFunction_STATE3[133]), .B(
        RoundFunction_STATE3[173]), .ZN(RoundFunction_T3_n413) );
  XOR2_X1 RoundFunction_T3_U21 ( .A(RoundFunction_STATE3[13]), .B(
        RoundFunction_STATE3[93]), .Z(RoundFunction_T3_n414) );
  XNOR2_X1 RoundFunction_T3_U20 ( .A(RoundFunction_STATE3[100]), .B(
        RoundFunction_T3_n561), .ZN(RoundFunction_TMP3_3[23]) );
  XNOR2_X1 RoundFunction_T3_U19 ( .A(RoundFunction_T3_n536), .B(
        RoundFunction_T3_n498), .ZN(RoundFunction_T3_n561) );
  XOR2_X1 RoundFunction_T3_U18 ( .A(RoundFunction_STATE3[107]), .B(
        RoundFunction_T3_n412), .Z(RoundFunction_T3_n498) );
  XNOR2_X1 RoundFunction_T3_U17 ( .A(RoundFunction_T3_n411), .B(
        RoundFunction_T3_n410), .ZN(RoundFunction_T3_n412) );
  XNOR2_X1 RoundFunction_T3_U16 ( .A(RoundFunction_STATE3[187]), .B(
        RoundFunction_STATE3[67]), .ZN(RoundFunction_T3_n410) );
  XOR2_X1 RoundFunction_T3_U15 ( .A(RoundFunction_STATE3[27]), .B(
        RoundFunction_STATE3[147]), .Z(RoundFunction_T3_n411) );
  XOR2_X1 RoundFunction_T3_U14 ( .A(RoundFunction_STATE3[52]), .B(
        RoundFunction_T3_n409), .Z(RoundFunction_T3_n536) );
  XNOR2_X1 RoundFunction_T3_U13 ( .A(RoundFunction_T3_n408), .B(
        RoundFunction_T3_n407), .ZN(RoundFunction_T3_n409) );
  XNOR2_X1 RoundFunction_T3_U12 ( .A(RoundFunction_STATE3[12]), .B(
        RoundFunction_STATE3[172]), .ZN(RoundFunction_T3_n407) );
  XOR2_X1 RoundFunction_T3_U11 ( .A(RoundFunction_STATE3[132]), .B(
        RoundFunction_STATE3[92]), .Z(RoundFunction_T3_n408) );
  XNOR2_X1 RoundFunction_T3_U10 ( .A(RoundFunction_STATE3[0]), .B(
        RoundFunction_T3_n581), .ZN(RoundFunction_TMP3_3[0]) );
  XNOR2_X1 RoundFunction_T3_U9 ( .A(RoundFunction_T3_n438), .B(
        RoundFunction_T3_n428), .ZN(RoundFunction_T3_n581) );
  XOR2_X1 RoundFunction_T3_U8 ( .A(RoundFunction_STATE3[55]), .B(
        RoundFunction_T3_n406), .Z(RoundFunction_T3_n428) );
  XNOR2_X1 RoundFunction_T3_U7 ( .A(RoundFunction_T3_n405), .B(
        RoundFunction_T3_n404), .ZN(RoundFunction_T3_n406) );
  XNOR2_X1 RoundFunction_T3_U6 ( .A(RoundFunction_STATE3[135]), .B(
        RoundFunction_STATE3[175]), .ZN(RoundFunction_T3_n404) );
  XOR2_X1 RoundFunction_T3_U5 ( .A(RoundFunction_STATE3[15]), .B(
        RoundFunction_STATE3[95]), .Z(RoundFunction_T3_n405) );
  XOR2_X1 RoundFunction_T3_U4 ( .A(RoundFunction_STATE3[112]), .B(
        RoundFunction_T3_n403), .Z(RoundFunction_T3_n438) );
  XNOR2_X1 RoundFunction_T3_U3 ( .A(RoundFunction_T3_n402), .B(
        RoundFunction_T3_n401), .ZN(RoundFunction_T3_n403) );
  XNOR2_X1 RoundFunction_T3_U2 ( .A(RoundFunction_STATE3[192]), .B(
        RoundFunction_STATE3[72]), .ZN(RoundFunction_T3_n401) );
  XOR2_X1 RoundFunction_T3_U1 ( .A(RoundFunction_STATE3[32]), .B(
        RoundFunction_STATE3[152]), .Z(RoundFunction_T3_n402) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_0_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_0_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[2]), .ZN(RESULT1[160]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[5]), .ZN(RESULT2[160]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[8]), .ZN(RESULT3[160]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[11]), .ZN(RESULT1[168]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[14]), .ZN(RESULT2[168]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[17]), .ZN(RESULT3[168]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[20]), .ZN(RESULT1[176]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[23]), .ZN(RESULT2[176]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[26]), .ZN(RESULT3[176]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[29]), .ZN(RESULT1[184]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[32]), .ZN(RESULT2[184]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[35]), .ZN(RESULT3[184]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[38]), .ZN(
        RoundFunction_TMP4_1[0]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[41]), .ZN(RESULT2[192]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[44]), .ZN(RESULT3[192]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_0_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_0_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_1_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_1_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[2]), .ZN(RESULT1[161]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[5]), .ZN(RESULT2[161]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[8]), .ZN(RESULT3[161]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[11]), .ZN(RESULT1[169]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[14]), .ZN(RESULT2[169]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[17]), .ZN(RESULT3[169]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[20]), .ZN(RESULT1[177]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[23]), .ZN(RESULT2[177]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[26]), .ZN(RESULT3[177]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[29]), .ZN(RESULT1[185]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[32]), .ZN(RESULT2[185]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[35]), .ZN(RESULT3[185]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[38]), .ZN(
        RoundFunction_TMP4_1[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[41]), .ZN(RESULT2[193]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[44]), .ZN(RESULT3[193]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_1_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_1_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_2_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_2_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[2]), .ZN(RESULT1[162]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[5]), .ZN(RESULT2[162]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[8]), .ZN(RESULT3[162]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[11]), .ZN(RESULT1[170]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[14]), .ZN(RESULT2[170]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[17]), .ZN(RESULT3[170]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[20]), .ZN(RESULT1[178]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[23]), .ZN(RESULT2[178]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[26]), .ZN(RESULT3[178]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[29]), .ZN(RESULT1[186]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[32]), .ZN(RESULT2[186]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[35]), .ZN(RESULT3[186]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[38]), .ZN(
        RoundFunction_TMP4_1[2]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[41]), .ZN(RESULT2[194]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[44]), .ZN(RESULT3[194]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_2_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_2_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_3_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_3_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[2]), .ZN(RESULT1[163]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[5]), .ZN(RESULT2[163]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[8]), .ZN(RESULT3[163]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[11]), .ZN(RESULT1[171]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[14]), .ZN(RESULT2[171]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[17]), .ZN(RESULT3[171]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[20]), .ZN(RESULT1[179]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[23]), .ZN(RESULT2[179]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[26]), .ZN(RESULT3[179]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[29]), .ZN(RESULT1[187]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[32]), .ZN(RESULT2[187]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[35]), .ZN(RESULT3[187]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[38]), .ZN(
        RoundFunction_TMP4_1[3]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[41]), .ZN(RESULT2[195]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[44]), .ZN(RESULT3[195]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_3_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_3_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_4_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_4_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[2]), .ZN(RESULT1[164]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[5]), .ZN(RESULT2[164]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[8]), .ZN(RESULT3[164]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[11]), .ZN(RESULT1[172]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[14]), .ZN(RESULT2[172]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[17]), .ZN(RESULT3[172]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[20]), .ZN(RESULT1[180]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[23]), .ZN(RESULT2[180]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[26]), .ZN(RESULT3[180]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[29]), .ZN(RESULT1[188]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[32]), .ZN(RESULT2[188]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[35]), .ZN(RESULT3[188]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[38]), .ZN(
        RoundFunction_TMP4_1[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[41]), .ZN(RESULT2[196]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[44]), .ZN(RESULT3[196]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_4_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_4_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_5_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_5_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[2]), .ZN(RESULT1[165]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[5]), .ZN(RESULT2[165]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[8]), .ZN(RESULT3[165]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[11]), .ZN(RESULT1[173]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[14]), .ZN(RESULT2[173]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[17]), .ZN(RESULT3[173]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[20]), .ZN(RESULT1[181]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[23]), .ZN(RESULT2[181]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[26]), .ZN(RESULT3[181]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[29]), .ZN(RESULT1[189]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[32]), .ZN(RESULT2[189]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[35]), .ZN(RESULT3[189]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[38]), .ZN(
        RoundFunction_TMP4_1[5]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[41]), .ZN(RESULT2[197]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[44]), .ZN(RESULT3[197]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_5_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_5_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_6_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_6_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[2]), .ZN(RESULT1[166]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[5]), .ZN(RESULT2[166]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[8]), .ZN(RESULT3[166]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[11]), .ZN(RESULT1[174]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[14]), .ZN(RESULT2[174]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[17]), .ZN(RESULT3[174]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[20]), .ZN(RESULT1[182]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[23]), .ZN(RESULT2[182]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[26]), .ZN(RESULT3[182]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[29]), .ZN(RESULT1[190]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[32]), .ZN(RESULT2[190]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[35]), .ZN(RESULT3[190]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[38]), .ZN(
        RoundFunction_TMP4_1[6]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[41]), .ZN(RESULT2[198]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[44]), .ZN(RESULT3[198]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_6_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_6_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_7_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_7_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[2]), .ZN(RESULT1[167]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[5]), .ZN(RESULT2[167]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[8]), .ZN(RESULT3[167]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[11]), .ZN(RESULT1[175]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[14]), .ZN(RESULT2[175]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[17]), .ZN(RESULT3[175]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[20]), .ZN(RESULT1[183]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[23]), .ZN(RESULT2[183]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[26]), .ZN(RESULT3[183]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[29]), .ZN(RESULT1[191]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[32]), .ZN(RESULT2[191]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[35]), .ZN(RESULT3[191]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[38]), .ZN(
        RoundFunction_TMP4_1[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[41]), .ZN(RESULT2[199]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[44]), .ZN(RESULT3[199]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_7_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_7_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[64]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[48]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[56]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[72]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[72]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[48]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[56]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[56]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[48]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[64]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[64]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[72]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_8_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_8_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[2]), .ZN(RESULT1[120]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[5]), .ZN(RESULT2[120]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[8]), .ZN(RESULT3[120]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[11]), .ZN(RESULT1[128]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[14]), .ZN(RESULT2[128]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[17]), .ZN(RESULT3[128]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[20]), .ZN(RESULT1[136]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[23]), .ZN(RESULT2[136]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[26]), .ZN(RESULT3[136]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[29]), .ZN(RESULT1[144]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[32]), .ZN(RESULT2[144]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[35]), .ZN(RESULT3[144]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[38]), .ZN(RESULT1[152]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[41]), .ZN(RESULT2[152]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[44]), .ZN(RESULT3[152]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_8_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_8_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[65]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[49]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[57]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[73]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[73]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[49]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[57]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[57]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[49]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[65]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[65]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[73]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_9_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_9_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[2]), .ZN(RESULT1[121]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[5]), .ZN(RESULT2[121]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[8]), .ZN(RESULT3[121]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[11]), .ZN(RESULT1[129]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[14]), .ZN(RESULT2[129]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[17]), .ZN(RESULT3[129]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[20]), .ZN(RESULT1[137]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[23]), .ZN(RESULT2[137]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[26]), .ZN(RESULT3[137]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[29]), .ZN(RESULT1[145]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[32]), .ZN(RESULT2[145]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[35]), .ZN(RESULT3[145]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression1_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression1_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[38]), .ZN(RESULT1[153]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression1_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression2_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression2_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[41]), .ZN(RESULT2[153]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression2_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression3_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression3_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[44]), .ZN(RESULT3[153]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression3_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_9_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_9_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[66]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[50]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[58]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[74]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[74]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[50]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[58]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[58]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[50]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[66]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[66]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[74]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_10_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_10_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_10_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[2]), .ZN(RESULT1[122])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[5]), .ZN(RESULT2[122])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[8]), .ZN(RESULT3[122])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[11]), .ZN(RESULT1[130])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[14]), .ZN(RESULT2[130])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[17]), .ZN(RESULT3[130])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[20]), .ZN(RESULT1[138])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[23]), .ZN(RESULT2[138])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[26]), .ZN(RESULT3[138])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[29]), .ZN(RESULT1[146])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[32]), .ZN(RESULT2[146])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[35]), .ZN(RESULT3[146])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[38]), .ZN(RESULT1[154])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[41]), .ZN(RESULT2[154])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[44]), .ZN(RESULT3[154])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_10_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_10_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[67]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[51]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[59]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[75]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[75]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[51]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[59]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[59]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[51]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[67]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[67]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[75]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_11_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_11_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_11_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[2]), .ZN(RESULT1[123])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[5]), .ZN(RESULT2[123])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[8]), .ZN(RESULT3[123])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[11]), .ZN(RESULT1[131])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[14]), .ZN(RESULT2[131])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[17]), .ZN(RESULT3[131])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[20]), .ZN(RESULT1[139])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[23]), .ZN(RESULT2[139])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[26]), .ZN(RESULT3[139])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[29]), .ZN(RESULT1[147])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[32]), .ZN(RESULT2[147])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[35]), .ZN(RESULT3[147])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[38]), .ZN(RESULT1[155])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[41]), .ZN(RESULT2[155])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[44]), .ZN(RESULT3[155])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_11_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_11_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[68]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[52]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[60]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[76]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[76]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[52]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[60]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[60]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[52]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[68]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[68]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[76]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_12_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_12_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_12_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[2]), .ZN(RESULT1[124])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[5]), .ZN(RESULT2[124])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[8]), .ZN(RESULT3[124])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[11]), .ZN(RESULT1[132])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[14]), .ZN(RESULT2[132])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[17]), .ZN(RESULT3[132])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[20]), .ZN(RESULT1[140])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[23]), .ZN(RESULT2[140])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[26]), .ZN(RESULT3[140])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[29]), .ZN(RESULT1[148])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[32]), .ZN(RESULT2[148])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[35]), .ZN(RESULT3[148])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[38]), .ZN(RESULT1[156])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[41]), .ZN(RESULT2[156])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[44]), .ZN(RESULT3[156])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_12_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_12_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[69]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[45]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[53]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[61]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[77]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[77]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[53]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[61]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[61]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[45]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[53]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[45]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[69]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[69]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[77]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_13_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_13_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_13_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[2]), .ZN(RESULT1[125])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[5]), .ZN(RESULT2[125])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[8]), .ZN(RESULT3[125])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[11]), .ZN(RESULT1[133])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[14]), .ZN(RESULT2[133])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[17]), .ZN(RESULT3[133])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[20]), .ZN(RESULT1[141])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[23]), .ZN(RESULT2[141])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[26]), .ZN(RESULT3[141])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[29]), .ZN(RESULT1[149])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[32]), .ZN(RESULT2[149])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[35]), .ZN(RESULT3[149])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[38]), .ZN(RESULT1[157])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[41]), .ZN(RESULT2[157])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[44]), .ZN(RESULT3[157])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_13_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_13_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[70]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[46]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[54]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[62]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[78]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[78]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[54]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[62]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[62]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[46]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[54]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[46]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[70]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[70]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[78]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_14_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_14_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_14_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[2]), .ZN(RESULT1[126])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[5]), .ZN(RESULT2[126])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[8]), .ZN(RESULT3[126])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[11]), .ZN(RESULT1[134])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[14]), .ZN(RESULT2[134])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[17]), .ZN(RESULT3[134])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[20]), .ZN(RESULT1[142])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[23]), .ZN(RESULT2[142])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[26]), .ZN(RESULT3[142])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[29]), .ZN(RESULT1[150])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[32]), .ZN(RESULT2[150])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[35]), .ZN(RESULT3[150])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[38]), .ZN(RESULT1[158])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[41]), .ZN(RESULT2[158])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[44]), .ZN(RESULT3[158])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_14_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_14_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[71]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[47]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[55]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[63]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[79]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[79]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[55]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[63]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[63]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[47]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[55]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[47]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[71]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[71]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[79]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_15_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_15_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_15_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[2]), .ZN(RESULT1[127])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[5]), .ZN(RESULT2[127])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[8]), .ZN(RESULT3[127])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[11]), .ZN(RESULT1[135])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[14]), .ZN(RESULT2[135])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[17]), .ZN(RESULT3[135])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[20]), .ZN(RESULT1[143])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[23]), .ZN(RESULT2[143])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[26]), .ZN(RESULT3[143])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[29]), .ZN(RESULT1[151])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[32]), .ZN(RESULT2[151])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[35]), .ZN(RESULT3[151])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[38]), .ZN(RESULT1[159])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[41]), .ZN(RESULT2[159])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[44]), .ZN(RESULT3[159])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_15_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_15_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[104]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[80]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[88]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[96]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[112]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[112]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[88]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[96]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[96]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[80]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[88]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[80]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[104]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[104]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[112]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_16_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_16_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_16_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[2]), .ZN(RESULT1[80]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[5]), .ZN(RESULT2[80]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[8]), .ZN(RESULT3[80]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[11]), .ZN(RESULT1[88])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[14]), .ZN(RESULT2[88])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[17]), .ZN(RESULT3[88])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[20]), .ZN(RESULT1[96])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[23]), .ZN(RESULT2[96])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[26]), .ZN(RESULT3[96])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[29]), .ZN(RESULT1[104])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[32]), .ZN(RESULT2[104])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[35]), .ZN(RESULT3[104])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[38]), .ZN(RESULT1[112])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[41]), .ZN(RESULT2[112])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[44]), .ZN(RESULT3[112])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_16_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_16_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[105]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[81]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[89]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[97]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[113]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[113]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[89]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[97]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[97]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[81]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[89]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[81]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[105]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[105]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[113]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_17_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_17_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_17_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[2]), .ZN(RESULT1[81]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[5]), .ZN(RESULT2[81]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[8]), .ZN(RESULT3[81]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[11]), .ZN(RESULT1[89])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[14]), .ZN(RESULT2[89])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[17]), .ZN(RESULT3[89])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[20]), .ZN(RESULT1[97])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[23]), .ZN(RESULT2[97])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[26]), .ZN(RESULT3[97])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[29]), .ZN(RESULT1[105])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[32]), .ZN(RESULT2[105])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[35]), .ZN(RESULT3[105])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[38]), .ZN(RESULT1[113])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[41]), .ZN(RESULT2[113])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[44]), .ZN(RESULT3[113])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_17_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_17_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[106]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[82]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[90]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[98]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[114]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[114]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[90]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[98]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[98]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[82]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[90]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[82]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[106]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[106]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[114]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_18_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_18_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_18_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[2]), .ZN(RESULT1[82]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[5]), .ZN(RESULT2[82]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[8]), .ZN(RESULT3[82]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[11]), .ZN(RESULT1[90])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[14]), .ZN(RESULT2[90])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[17]), .ZN(RESULT3[90])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[20]), .ZN(RESULT1[98])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[23]), .ZN(RESULT2[98])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[26]), .ZN(RESULT3[98])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[29]), .ZN(RESULT1[106])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[32]), .ZN(RESULT2[106])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[35]), .ZN(RESULT3[106])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[38]), .ZN(RESULT1[114])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[41]), .ZN(RESULT2[114])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[44]), .ZN(RESULT3[114])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_18_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_18_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[107]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[83]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[91]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[99]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[115]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[115]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[91]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[99]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[99]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[83]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[91]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[83]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[107]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[107]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[115]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_19_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_19_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_19_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[2]), .ZN(RESULT1[83]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[5]), .ZN(RESULT2[83]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[8]), .ZN(RESULT3[83]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[11]), .ZN(RESULT1[91])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[14]), .ZN(RESULT2[91])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[17]), .ZN(RESULT3[91])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[20]), .ZN(RESULT1[99])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[23]), .ZN(RESULT2[99])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[26]), .ZN(RESULT3[99])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[29]), .ZN(RESULT1[107])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[32]), .ZN(RESULT2[107])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[35]), .ZN(RESULT3[107])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[38]), .ZN(RESULT1[115])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[41]), .ZN(RESULT2[115])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[44]), .ZN(RESULT3[115])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_19_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_19_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[108]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[84]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[92]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[100]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[116]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[116]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[92]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[100]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[100]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[84]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[92]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[84]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[108]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[108]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[116]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_20_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_20_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_20_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[2]), .ZN(RESULT1[84]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[5]), .ZN(RESULT2[84]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[8]), .ZN(RESULT3[84]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[11]), .ZN(RESULT1[92])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[14]), .ZN(RESULT2[92])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[17]), .ZN(RESULT3[92])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[20]), .ZN(RESULT1[100])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[23]), .ZN(RESULT2[100])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[26]), .ZN(RESULT3[100])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[29]), .ZN(RESULT1[108])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[32]), .ZN(RESULT2[108])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[35]), .ZN(RESULT3[108])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[38]), .ZN(RESULT1[116])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[41]), .ZN(RESULT2[116])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[44]), .ZN(RESULT3[116])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_20_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_20_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[109]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[85]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[93]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[101]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[117]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[117]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[93]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[101]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[101]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[85]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[93]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[85]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[109]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[109]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[117]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_21_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_21_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_21_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[2]), .ZN(RESULT1[85]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[5]), .ZN(RESULT2[85]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[8]), .ZN(RESULT3[85]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[11]), .ZN(RESULT1[93])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[14]), .ZN(RESULT2[93])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[17]), .ZN(RESULT3[93])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[20]), .ZN(RESULT1[101])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[23]), .ZN(RESULT2[101])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[26]), .ZN(RESULT3[101])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[29]), .ZN(RESULT1[109])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[32]), .ZN(RESULT2[109])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[35]), .ZN(RESULT3[109])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[38]), .ZN(RESULT1[117])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[41]), .ZN(RESULT2[117])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[44]), .ZN(RESULT3[117])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_21_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_21_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[110]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[86]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[94]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[102]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[118]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[118]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[94]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[102]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[102]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[86]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[94]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[86]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[110]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[110]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[118]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_22_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_22_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_22_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[2]), .ZN(RESULT1[86]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[5]), .ZN(RESULT2[86]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[8]), .ZN(RESULT3[86]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[11]), .ZN(RESULT1[94])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[14]), .ZN(RESULT2[94])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[17]), .ZN(RESULT3[94])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[20]), .ZN(RESULT1[102])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[23]), .ZN(RESULT2[102])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[26]), .ZN(RESULT3[102])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[29]), .ZN(RESULT1[110])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[32]), .ZN(RESULT2[110])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[35]), .ZN(RESULT3[110])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[38]), .ZN(RESULT1[118])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[41]), .ZN(RESULT2[118])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[44]), .ZN(RESULT3[118])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_22_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_22_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[111]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[87]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[95]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[103]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[119]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[119]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[95]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[103]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[103]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[87]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[95]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[87]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[111]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[111]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[119]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_23_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_23_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_23_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[2]), .ZN(RESULT1[87]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[5]), .ZN(RESULT2[87]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[8]), .ZN(RESULT3[87]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[11]), .ZN(RESULT1[95])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[14]), .ZN(RESULT2[95])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[17]), .ZN(RESULT3[95])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[20]), .ZN(RESULT1[103])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[23]), .ZN(RESULT2[103])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[26]), .ZN(RESULT3[103])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[29]), .ZN(RESULT1[111])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[32]), .ZN(RESULT2[111])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[35]), .ZN(RESULT3[111])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[38]), .ZN(RESULT1[119])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[41]), .ZN(RESULT2[119])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[44]), .ZN(RESULT3[119])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_23_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_23_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[144]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[120]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[128]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[136]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[152]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[152]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[128]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[136]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[136]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[120]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[128]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[120]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[144]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[144]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[152]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_24_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_24_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_24_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[2]), .ZN(RESULT1[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[5]), .ZN(RESULT2[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[8]), .ZN(RESULT3[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[11]), .ZN(RESULT1[48])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[14]), .ZN(RESULT2[48])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[17]), .ZN(RESULT3[48])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[20]), .ZN(RESULT1[56])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[23]), .ZN(RESULT2[56])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[26]), .ZN(RESULT3[56])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[29]), .ZN(RESULT1[64])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[32]), .ZN(RESULT2[64])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[35]), .ZN(RESULT3[64])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[38]), .ZN(RESULT1[72])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[41]), .ZN(RESULT2[72])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[44]), .ZN(RESULT3[72])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_24_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_24_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[145]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[121]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[129]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[137]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[153]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[153]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[129]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[137]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[137]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[121]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[129]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[121]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[145]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[145]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[153]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_25_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_25_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_25_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[2]), .ZN(RESULT1[41]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[5]), .ZN(RESULT2[41]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[8]), .ZN(RESULT3[41]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[11]), .ZN(RESULT1[49])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[14]), .ZN(RESULT2[49])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[17]), .ZN(RESULT3[49])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[20]), .ZN(RESULT1[57])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[23]), .ZN(RESULT2[57])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[26]), .ZN(RESULT3[57])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[29]), .ZN(RESULT1[65])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[32]), .ZN(RESULT2[65])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[35]), .ZN(RESULT3[65])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[38]), .ZN(RESULT1[73])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[41]), .ZN(RESULT2[73])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[44]), .ZN(RESULT3[73])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_25_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_25_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[146]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[122]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[130]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[138]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[154]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[154]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[130]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[138]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[138]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[122]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[130]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[122]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[146]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[146]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[154]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_26_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_26_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_26_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[2]), .ZN(RESULT1[42]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[5]), .ZN(RESULT2[42]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[8]), .ZN(RESULT3[42]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[11]), .ZN(RESULT1[50])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[14]), .ZN(RESULT2[50])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[17]), .ZN(RESULT3[50])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[20]), .ZN(RESULT1[58])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[23]), .ZN(RESULT2[58])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[26]), .ZN(RESULT3[58])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[29]), .ZN(RESULT1[66])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[32]), .ZN(RESULT2[66])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[35]), .ZN(RESULT3[66])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[38]), .ZN(RESULT1[74])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[41]), .ZN(RESULT2[74])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[44]), .ZN(RESULT3[74])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_26_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_26_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[147]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[123]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[131]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[139]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[155]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[155]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[131]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[139]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[139]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[123]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[131]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[123]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[147]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[147]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[155]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_27_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_27_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_27_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[2]), .ZN(RESULT1[43]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[5]), .ZN(RESULT2[43]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[8]), .ZN(RESULT3[43]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[11]), .ZN(RESULT1[51])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[14]), .ZN(RESULT2[51])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[17]), .ZN(RESULT3[51])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[20]), .ZN(RESULT1[59])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[23]), .ZN(RESULT2[59])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[26]), .ZN(RESULT3[59])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[29]), .ZN(RESULT1[67])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[32]), .ZN(RESULT2[67])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[35]), .ZN(RESULT3[67])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[38]), .ZN(RESULT1[75])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[41]), .ZN(RESULT2[75])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[44]), .ZN(RESULT3[75])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_27_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_27_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[148]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[124]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[132]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[140]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[156]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[156]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[132]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[140]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[140]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[124]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[132]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[124]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[148]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[148]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[156]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_28_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_28_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_28_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[2]), .ZN(RESULT1[44]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[5]), .ZN(RESULT2[44]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[8]), .ZN(RESULT3[44]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[11]), .ZN(RESULT1[52])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[14]), .ZN(RESULT2[52])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[17]), .ZN(RESULT3[52])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[20]), .ZN(RESULT1[60])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[23]), .ZN(RESULT2[60])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[26]), .ZN(RESULT3[60])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[29]), .ZN(RESULT1[68])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[32]), .ZN(RESULT2[68])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[35]), .ZN(RESULT3[68])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[38]), .ZN(RESULT1[76])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[41]), .ZN(RESULT2[76])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[44]), .ZN(RESULT3[76])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_28_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_28_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[149]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[125]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[133]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[141]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[157]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[157]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[133]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[141]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[141]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[125]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[133]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[125]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[149]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[149]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[157]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_29_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_29_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_29_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[2]), .ZN(RESULT1[45]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[5]), .ZN(RESULT2[45]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[8]), .ZN(RESULT3[45]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[11]), .ZN(RESULT1[53])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[14]), .ZN(RESULT2[53])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[17]), .ZN(RESULT3[53])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[20]), .ZN(RESULT1[61])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[23]), .ZN(RESULT2[61])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[26]), .ZN(RESULT3[61])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[29]), .ZN(RESULT1[69])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[32]), .ZN(RESULT2[69])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[35]), .ZN(RESULT3[69])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[38]), .ZN(RESULT1[77])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[41]), .ZN(RESULT2[77])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[44]), .ZN(RESULT3[77])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_29_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_29_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[150]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[126]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[134]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[142]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[158]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[158]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[134]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[142]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[142]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[126]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[134]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[126]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[150]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[150]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[158]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_30_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_30_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_30_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[2]), .ZN(RESULT1[46]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[5]), .ZN(RESULT2[46]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[8]), .ZN(RESULT3[46]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[11]), .ZN(RESULT1[54])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[14]), .ZN(RESULT2[54])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[17]), .ZN(RESULT3[54])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[20]), .ZN(RESULT1[62])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[23]), .ZN(RESULT2[62])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[26]), .ZN(RESULT3[62])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[29]), .ZN(RESULT1[70])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[32]), .ZN(RESULT2[70])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[35]), .ZN(RESULT3[70])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[38]), .ZN(RESULT1[78])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[41]), .ZN(RESULT2[78])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[44]), .ZN(RESULT3[78])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_30_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_30_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[151]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[127]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[135]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[143]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[159]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[159]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[135]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[143]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[143]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[127]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[135]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[127]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[151]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[151]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[159]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_31_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_31_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_31_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[2]), .ZN(RESULT1[47]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[5]), .ZN(RESULT2[47]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[8]), .ZN(RESULT3[47]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[11]), .ZN(RESULT1[55])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[14]), .ZN(RESULT2[55])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[17]), .ZN(RESULT3[55])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[20]), .ZN(RESULT1[63])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[23]), .ZN(RESULT2[63])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[26]), .ZN(RESULT3[63])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[29]), .ZN(RESULT1[71])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[32]), .ZN(RESULT2[71])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[35]), .ZN(RESULT3[71])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[38]), .ZN(RESULT1[79])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[41]), .ZN(RESULT2[79])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[44]), .ZN(RESULT3[79])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_31_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_31_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[184]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[160]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[168]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[176]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[192]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[192]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[168]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[176]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[176]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[160]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[168]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[160]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[184]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[184]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[192]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_32_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_32_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_32_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[2]), .ZN(RESULT1[0]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[5]), .ZN(RESULT2[0]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[8]), .ZN(RESULT3[0]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[11]), .ZN(RESULT1[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[14]), .ZN(RESULT2[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[17]), .ZN(RESULT3[8]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[20]), .ZN(RESULT1[16])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[23]), .ZN(RESULT2[16])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[26]), .ZN(RESULT3[16])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[29]), .ZN(RESULT1[24])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[32]), .ZN(RESULT2[24])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[35]), .ZN(RESULT3[24])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[38]), .ZN(RESULT1[32])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[41]), .ZN(RESULT2[32])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[44]), .ZN(RESULT3[32])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_32_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_32_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[185]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[161]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[169]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[177]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[193]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[193]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[169]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[177]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[177]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[161]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[169]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[161]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[185]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[185]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[193]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_33_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_33_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_33_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[2]), .ZN(RESULT1[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[5]), .ZN(RESULT2[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[8]), .ZN(RESULT3[1]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[11]), .ZN(RESULT1[9]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[14]), .ZN(RESULT2[9]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[17]), .ZN(RESULT3[9]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[20]), .ZN(RESULT1[17])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[23]), .ZN(RESULT2[17])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[26]), .ZN(RESULT3[17])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[29]), .ZN(RESULT1[25])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[32]), .ZN(RESULT2[25])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[35]), .ZN(RESULT3[25])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[38]), .ZN(RESULT1[33])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[41]), .ZN(RESULT2[33])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[44]), .ZN(RESULT3[33])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_33_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_33_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[186]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[162]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[170]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[178]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[194]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[194]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[170]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[178]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[178]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[162]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[170]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[162]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[186]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[186]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[194]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_34_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_34_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_34_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[2]), .ZN(RESULT1[2]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[5]), .ZN(RESULT2[2]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[8]), .ZN(RESULT3[2]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[11]), .ZN(RESULT1[10])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[14]), .ZN(RESULT2[10])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[17]), .ZN(RESULT3[10])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[20]), .ZN(RESULT1[18])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[23]), .ZN(RESULT2[18])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[26]), .ZN(RESULT3[18])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[29]), .ZN(RESULT1[26])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[32]), .ZN(RESULT2[26])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[35]), .ZN(RESULT3[26])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[38]), .ZN(RESULT1[34])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[41]), .ZN(RESULT2[34])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[44]), .ZN(RESULT3[34])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_34_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_34_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[187]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[163]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[171]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[179]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[195]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[195]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[171]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[179]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[179]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[163]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[171]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[163]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[187]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[187]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[195]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_35_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_35_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_35_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[2]), .ZN(RESULT1[3]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[5]), .ZN(RESULT2[3]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[8]), .ZN(RESULT3[3]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[11]), .ZN(RESULT1[11])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[14]), .ZN(RESULT2[11])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[17]), .ZN(RESULT3[11])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[20]), .ZN(RESULT1[19])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[23]), .ZN(RESULT2[19])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[26]), .ZN(RESULT3[19])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[29]), .ZN(RESULT1[27])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[32]), .ZN(RESULT2[27])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[35]), .ZN(RESULT3[27])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[38]), .ZN(RESULT1[35])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[41]), .ZN(RESULT2[35])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[44]), .ZN(RESULT3[35])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_35_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_35_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[188]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[164]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[172]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[180]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[196]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[196]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[172]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[180]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[180]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[164]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[172]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[164]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[188]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[188]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[196]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_36_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_36_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_36_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[2]), .ZN(RESULT1[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[5]), .ZN(RESULT2[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[8]), .ZN(RESULT3[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[11]), .ZN(RESULT1[12])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[14]), .ZN(RESULT2[12])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[17]), .ZN(RESULT3[12])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[20]), .ZN(RESULT1[20])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[23]), .ZN(RESULT2[20])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[26]), .ZN(RESULT3[20])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[29]), .ZN(RESULT1[28])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[32]), .ZN(RESULT2[28])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[35]), .ZN(RESULT3[28])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[38]), .ZN(RESULT1[36])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[41]), .ZN(RESULT2[36])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[44]), .ZN(RESULT3[36])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_36_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_36_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[189]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[165]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[173]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[181]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[197]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[197]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[173]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[181]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[181]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[165]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[173]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[165]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[189]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[189]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[197]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_37_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_37_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_37_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[2]), .ZN(RESULT1[5]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[5]), .ZN(RESULT2[5]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[8]), .ZN(RESULT3[5]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[11]), .ZN(RESULT1[13])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[14]), .ZN(RESULT2[13])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[17]), .ZN(RESULT3[13])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[20]), .ZN(RESULT1[21])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[23]), .ZN(RESULT2[21])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[26]), .ZN(RESULT3[21])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[29]), .ZN(RESULT1[29])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[32]), .ZN(RESULT2[29])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[35]), .ZN(RESULT3[29])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[38]), .ZN(RESULT1[37])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[41]), .ZN(RESULT2[37])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[44]), .ZN(RESULT3[37])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_37_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_37_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[190]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[166]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[174]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[182]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[198]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[198]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[174]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[182]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[182]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[166]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[174]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[166]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[190]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[190]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[198]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_38_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_38_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_38_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[2]), .ZN(RESULT1[6]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[5]), .ZN(RESULT2[6]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[8]), .ZN(RESULT3[6]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[11]), .ZN(RESULT1[14])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[14]), .ZN(RESULT2[14])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[17]), .ZN(RESULT3[14])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[20]), .ZN(RESULT1[22])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[23]), .ZN(RESULT2[22])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[26]), .ZN(RESULT3[22])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[29]), .ZN(RESULT1[30])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[32]), .ZN(RESULT2[30])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[35]), .ZN(RESULT3[30])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[38]), .ZN(RESULT1[38])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[41]), .ZN(RESULT2[38])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[44]), .ZN(RESULT3[38])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_38_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_38_InstXOR_4__Compression3_n3) );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_b_reg_3_ ( .D(
        RoundFunction_TMP3_3[191]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_e_reg_3_ ( .D(
        RoundFunction_TMP3_3[167]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_d_reg_3_ ( .D(
        RoundFunction_TMP3_3[175]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_c_reg_3_ ( .D(
        RoundFunction_TMP3_3[183]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_a_reg_1_ ( .D(
        RoundFunction_TMP3_1[199]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_a_reg_2_ ( .D(
        RoundFunction_TMP3_2[199]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_d_reg_1_ ( .D(
        RoundFunction_TMP3_1[175]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_c_reg_1_ ( .D(
        RoundFunction_TMP3_1[183]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_c_reg_2_ ( .D(
        RoundFunction_TMP3_2[183]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_e_reg_2_ ( .D(
        RoundFunction_TMP3_2[167]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_d_reg_2_ ( .D(
        RoundFunction_TMP3_2[175]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_e_reg_1_ ( .D(
        RoundFunction_TMP3_1[167]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_b_reg_1_ ( .D(
        RoundFunction_TMP3_1[191]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_1_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_b_reg_2_ ( .D(
        RoundFunction_TMP3_2[191]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_2_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_a_reg_3_ ( .D(
        RoundFunction_TMP3_3[199]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_3_), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_0_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[0]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[0]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_1_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[1]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[1]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_2_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[2]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[2]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_3_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[3]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[3]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_4_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[4]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[4]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_5_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[5]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[5]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_6_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[6]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[6]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_7_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[7]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[7]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_8_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[8]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[8]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_9_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[9]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[9]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_10_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[10]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[10]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_11_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[11]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[11]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_12_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[12]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[12]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_13_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[13]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[13]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_14_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[14]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[14]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_15_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[15]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[15]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_16_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[16]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[16]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_17_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[17]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[17]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_18_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[18]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[18]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_19_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[19]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[19]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_20_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[20]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[20]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_21_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[21]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[21]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_22_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[22]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[22]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_23_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[23]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[23]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_24_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[24]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[24]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_25_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[25]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[25]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_26_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[26]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[26]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_27_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[27]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[27]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_28_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[28]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[28]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_29_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[29]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[29]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_30_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[30]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[30]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_31_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[31]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[31]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_32_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[32]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[32]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_33_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[33]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[33]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_34_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[34]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[34]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_35_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[35]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[35]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_36_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[36]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[36]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_37_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[37]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[37]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_38_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[38]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[38]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_39_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[39]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[39]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_40_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[40]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[40]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_41_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[41]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[41]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_42_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[42]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[42]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_43_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[43]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[43]), .QN() );
  DFF_X1 RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg_reg_44_ ( .D(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[44]), .CK(CLK), .Q(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[44]), .QN() );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[0]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_0__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_1__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_1__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[1]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_1__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_1__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_2__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[2]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_3__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_3__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[3]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_3__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_3__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_4__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[4]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_5__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_5__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[5]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_5__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_5__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_6__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_6__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[6]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_6__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_6__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_7__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_8__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_8__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[8]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_8__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_8__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_8__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_8__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_8__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_9__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_9__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[9]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_9__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_9__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_10__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_10__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[10]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_10__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_10__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_11__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_11__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[11]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_11__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_11__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_12__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_12__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[12]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_12__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_12__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_13__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[13]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_14__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_14__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[14]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_14__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_14__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_14__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_14__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_14__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_15__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_15__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[15]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_15__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_15__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_16__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[16]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_17__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_17__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[17]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_17__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_17__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[18]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_18__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[19]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_19__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_20__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_20__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[20]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_20__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_20__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_21__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_21__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[21]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_21__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_21__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_22__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[22]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_23__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_23__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[23]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_23__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_23__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_24__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_24__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[24]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_24__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_24__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_24__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_24__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_24__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_25__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_25__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[25]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_25__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_25__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_26__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_a_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[26]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_27__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[27]) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_28__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[28]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_29__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_3_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_29__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[29]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_29__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_29__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_29__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_29__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_29__CF_Inst_n5) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_30__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_30__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[30]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_30__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_30__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_31__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[31]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_32__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_1_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_32__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[32]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_32__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_32__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_32__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_32__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_32__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_33__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_33__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[33]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_33__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_33__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_34__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_34__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[34]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_34__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_34__CF_Inst_n3) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_35__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_b_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_35__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[35]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_35__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_35__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_36__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[36]) );
  OR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_37__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[37]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_38__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_38__CF_Inst_n7), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[38]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_38__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_38__CF_Inst_n7) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_39__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_39__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[39]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_39__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_1_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_39__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_40__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[40]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_41__CF_Inst_U3 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_2_), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_41__CF_Inst_n6), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[41]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_41__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_41__CF_Inst_n5), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_41__CF_Inst_n6) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_41__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_2_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_41__CF_Inst_n5) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_42__CF_Inst_U2 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_42__CF_Inst_n3), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_e_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[42]) );
  NAND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_42__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_1_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_42__CF_Inst_n3) );
  AND2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_43__CF_Inst_U1 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_2_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[43]) );
  NOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_44__CF_Inst_U2 ( .A1(
        RoundFunction_C_Inst_Chi_NoFresh_39_d_3_), .A2(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_44__CF_Inst_n3), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Out[44]) );
  INV_X1 RoundFunction_C_Inst_Chi_NoFresh_39_Inst_44__CF_Inst_U1 ( .A(
        RoundFunction_C_Inst_Chi_NoFresh_39_c_3_), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_Inst_44__CF_Inst_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[2]), .ZN(RESULT1[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[0]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[1]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[5]), .ZN(RESULT2[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[3]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[4]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[8]), .ZN(RESULT3[7]) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[6]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[7]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_0__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[11]), .ZN(RESULT1[15])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[9]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[10]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[14]), .ZN(RESULT2[15])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[12]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[13]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[17]), .ZN(RESULT3[15])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[15]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[16]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_1__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[20]), .ZN(RESULT1[23])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[18]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[19]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[23]), .ZN(RESULT2[23])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[21]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[22]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[26]), .ZN(RESULT3[23])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[24]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[25]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_2__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[29]), .ZN(RESULT1[31])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[27]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[28]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[32]), .ZN(RESULT2[31])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[30]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[31]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[35]), .ZN(RESULT3[31])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[33]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[34]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_3__Compression3_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression1_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression1_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[38]), .ZN(RESULT1[39])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression1_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[36]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[37]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression1_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression2_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression2_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[41]), .ZN(RESULT2[39])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression2_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[39]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[40]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression2_n3) );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression3_U2 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression3_n3), 
        .B(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[44]), .ZN(RESULT3[39])
         );
  XNOR2_X1 RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression3_U1 ( 
        .A(RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[42]), .B(
        RoundFunction_C_Inst_Chi_NoFresh_39_CF_Reg[43]), .ZN(
        RoundFunction_C_Inst_Chi_NoFresh_39_InstXOR_4__Compression3_n3) );
  OAI22_X1 FSM_U71 ( .A1(RESET), .A2(FSM_n92), .B1(FSM_n91), .B2(FSM_n90), 
        .ZN(FSM_n1) );
  AND3_X1 FSM_U70 ( .A1(FSM_n89), .A2(FSM_n88), .A3(FSM_n91), .ZN(FSM_n79) );
  OR2_X1 FSM_U69 ( .A1(FSM_n86), .A2(FSM_n85), .ZN(FSM_n91) );
  AOI221_X1 FSM_U68 ( .B1(FSM_n84), .B2(FSM_n88), .C1(FSM_n85), .C2(FSM_n88), 
        .A(FSM_n90), .ZN(FSM_n78) );
  INV_X1 FSM_U67 ( .A(FSM_n89), .ZN(FSM_n90) );
  NOR2_X1 FSM_U66 ( .A1(RESET), .A2(FSM_n87), .ZN(FSM_n89) );
  OR2_X1 FSM_U65 ( .A1(FSM_n28), .A2(FSM_n17), .ZN(FSM_n85) );
  INV_X1 FSM_U64 ( .A(FSM_n86), .ZN(FSM_n84) );
  OAI22_X1 FSM_U63 ( .A1(FSM_n8), .A2(FSM_n83), .B1(FSM_n7), .B2(FSM_n82), 
        .ZN(FSM_n77) );
  OAI221_X1 FSM_U62 ( .B1(FSM_n81), .B2(FSM_n80), .C1(FSM_n82), .C2(FSM_n15), 
        .A(FSM_n29), .ZN(FSM_n76) );
  XNOR2_X1 FSM_U61 ( .A(FSM_n69), .B(FSM_n68), .ZN(FSM_n80) );
  AOI22_X1 FSM_U60 ( .A1(FSM_n11), .A2(FSM_n12), .B1(FSM_n20), .B2(FSM_n22), 
        .ZN(FSM_n68) );
  OAI21_X1 FSM_U59 ( .B1(FSM_n10), .B2(FSM_n26), .A(FSM_n67), .ZN(FSM_n69) );
  INV_X1 FSM_U58 ( .A(FSM_n82), .ZN(FSM_n81) );
  OAI22_X1 FSM_U57 ( .A1(FSM_n15), .A2(FSM_n83), .B1(FSM_n14), .B2(FSM_n82), 
        .ZN(FSM_n75) );
  OAI22_X1 FSM_U56 ( .A1(FSM_n13), .A2(FSM_n82), .B1(FSM_n14), .B2(FSM_n83), 
        .ZN(FSM_n74) );
  OAI22_X1 FSM_U55 ( .A1(FSM_n12), .A2(FSM_n82), .B1(FSM_n13), .B2(FSM_n83), 
        .ZN(FSM_n73) );
  OAI22_X1 FSM_U54 ( .A1(FSM_n12), .A2(FSM_n83), .B1(FSM_n11), .B2(FSM_n82), 
        .ZN(FSM_n72) );
  OAI22_X1 FSM_U53 ( .A1(FSM_n10), .A2(FSM_n82), .B1(FSM_n11), .B2(FSM_n83), 
        .ZN(FSM_n71) );
  OAI22_X1 FSM_U52 ( .A1(FSM_n10), .A2(FSM_n83), .B1(FSM_n8), .B2(FSM_n82), 
        .ZN(FSM_n70) );
  NAND2_X1 FSM_U51 ( .A1(FSM_n29), .A2(FSM_n82), .ZN(FSM_n83) );
  NAND2_X1 FSM_U50 ( .A1(FSM_n17), .A2(FSM_n28), .ZN(FSM_n88) );
  INV_X1 FSM_U49 ( .A(FSM_n92), .ZN(DONE) );
  NAND3_X1 FSM_U48 ( .A1(FSM_n87), .A2(FSM_n17), .A3(FSM_n18), .ZN(FSM_n92) );
  NAND4_X1 FSM_U47 ( .A1(FSM_n66), .A2(FSM_n65), .A3(FSM_n64), .A4(FSM_n86), 
        .ZN(FSM_CONST_internal_7) );
  AOI21_X1 FSM_U46 ( .B1(FSM_n63), .B2(FSM_n62), .A(FSM_n61), .ZN(FSM_n65) );
  NOR3_X1 FSM_U45 ( .A1(FSM_n15), .A2(FSM_n11), .A3(FSM_n20), .ZN(FSM_n62) );
  NAND3_X1 FSM_U44 ( .A1(FSM_n60), .A2(FSM_n59), .A3(FSM_n64), .ZN(
        FSM_CONST_internal_3) );
  NAND3_X1 FSM_U43 ( .A1(FSM_n58), .A2(FSM_n57), .A3(FSM_n56), .ZN(FSM_n64) );
  NOR2_X1 FSM_U42 ( .A1(FSM_n55), .A2(FSM_n54), .ZN(FSM_n60) );
  NAND4_X1 FSM_U41 ( .A1(FSM_n66), .A2(FSM_n53), .A3(FSM_n59), .A4(FSM_n52), 
        .ZN(FSM_CONST_internal[1]) );
  NAND4_X1 FSM_U40 ( .A1(FSM_n13), .A2(FSM_n51), .A3(FSM_n20), .A4(FSM_n23), 
        .ZN(FSM_n52) );
  NAND4_X1 FSM_U39 ( .A1(FSM_n13), .A2(FSM_n15), .A3(FSM_n50), .A4(FSM_n49), 
        .ZN(FSM_n59) );
  NOR4_X1 FSM_U38 ( .A1(FSM_n14), .A2(FSM_n7), .A3(FSM_n10), .A4(FSM_n22), 
        .ZN(FSM_n49) );
  AOI21_X1 FSM_U37 ( .B1(FSM_n48), .B2(FSM_n47), .A(FSM_n55), .ZN(FSM_n66) );
  AOI221_X1 FSM_U36 ( .B1(FSM_n46), .B2(FSM_n45), .C1(FSM_n44), .C2(FSM_n45), 
        .A(FSM_n24), .ZN(FSM_n55) );
  AOI21_X1 FSM_U35 ( .B1(FSM_n10), .B2(FSM_n57), .A(FSM_n48), .ZN(FSM_n46) );
  NOR3_X1 FSM_U34 ( .A1(FSM_n11), .A2(FSM_n12), .A3(FSM_n43), .ZN(FSM_n57) );
  NAND2_X1 FSM_U33 ( .A1(FSM_n7), .A2(FSM_n8), .ZN(FSM_n43) );
  NOR2_X1 FSM_U32 ( .A1(FSM_n22), .A2(FSM_n42), .ZN(FSM_n48) );
  OR4_X1 FSM_U31 ( .A1(FSM_n41), .A2(FSM_n61), .A3(FSM_n54), .A4(FSM_n40), 
        .ZN(FSM_CONST_internal[0]) );
  OAI22_X1 FSM_U30 ( .A1(FSM_n45), .A2(FSM_n24), .B1(FSM_n56), .B2(FSM_n39), 
        .ZN(FSM_n40) );
  OAI211_X1 FSM_U29 ( .C1(FSM_n14), .C2(FSM_n27), .A(FSM_n13), .B(FSM_n38), 
        .ZN(FSM_n39) );
  AOI22_X1 FSM_U28 ( .A1(FSM_n37), .A2(FSM_n36), .B1(FSM_n35), .B2(FSM_n34), 
        .ZN(FSM_n45) );
  OAI33_X1 FSM_U27 ( .A1(FSM_n12), .A2(FSM_n33), .A3(FSM_n23), .B1(FSM_n20), 
        .B2(FSM_n44), .B3(FSM_n8), .ZN(FSM_n34) );
  NAND2_X1 FSM_U26 ( .A1(FSM_n15), .A2(FSM_n21), .ZN(FSM_n44) );
  NOR2_X1 FSM_U25 ( .A1(FSM_n22), .A2(FSM_n67), .ZN(FSM_n35) );
  INV_X1 FSM_U24 ( .A(FSM_n33), .ZN(FSM_n36) );
  OAI211_X1 FSM_U23 ( .C1(FSM_n33), .C2(FSM_n32), .A(FSM_n31), .B(FSM_n86), 
        .ZN(FSM_n54) );
  NAND2_X1 FSM_U22 ( .A1(FSM_n47), .A2(FSM_n37), .ZN(FSM_n86) );
  NOR2_X1 FSM_U21 ( .A1(FSM_n11), .A2(FSM_n42), .ZN(FSM_n37) );
  NAND4_X1 FSM_U20 ( .A1(FSM_n7), .A2(FSM_n8), .A3(FSM_n12), .A4(FSM_n10), 
        .ZN(FSM_n42) );
  AND2_X1 FSM_U19 ( .A1(FSM_n24), .A2(FSM_n58), .ZN(FSM_n47) );
  NOR2_X1 FSM_U18 ( .A1(FSM_n21), .A2(FSM_n25), .ZN(FSM_n58) );
  NAND4_X1 FSM_U17 ( .A1(FSM_n11), .A2(FSM_n15), .A3(FSM_n63), .A4(FSM_n20), 
        .ZN(FSM_n31) );
  NOR4_X1 FSM_U16 ( .A1(FSM_n14), .A2(FSM_n13), .A3(FSM_n23), .A4(FSM_n67), 
        .ZN(FSM_n63) );
  NAND2_X1 FSM_U15 ( .A1(FSM_n10), .A2(FSM_n26), .ZN(FSM_n67) );
  NAND4_X1 FSM_U14 ( .A1(FSM_n7), .A2(FSM_n50), .A3(FSM_n56), .A4(FSM_n22), 
        .ZN(FSM_n32) );
  NAND2_X1 FSM_U13 ( .A1(FSM_n25), .A2(FSM_n13), .ZN(FSM_n33) );
  AND3_X1 FSM_U12 ( .A1(FSM_n50), .A2(FSM_n51), .A3(FSM_n21), .ZN(FSM_n61) );
  NOR3_X1 FSM_U11 ( .A1(FSM_n14), .A2(FSM_n27), .A3(FSM_n30), .ZN(FSM_n51) );
  NOR2_X1 FSM_U10 ( .A1(FSM_n8), .A2(FSM_n20), .ZN(FSM_n50) );
  INV_X1 FSM_U9 ( .A(FSM_n53), .ZN(FSM_n41) );
  NAND3_X1 FSM_U8 ( .A1(FSM_n56), .A2(FSM_n38), .A3(FSM_n21), .ZN(FSM_n53) );
  NOR3_X1 FSM_U7 ( .A1(FSM_n23), .A2(FSM_n20), .A3(FSM_n30), .ZN(FSM_n38) );
  NAND3_X1 FSM_U6 ( .A1(FSM_n11), .A2(FSM_n7), .A3(FSM_n25), .ZN(FSM_n30) );
  NOR2_X1 FSM_U5 ( .A1(FSM_n10), .A2(FSM_n24), .ZN(FSM_n56) );
  INV_X1 FSM_U4 ( .A(RESET), .ZN(FSM_n29) );
  OAI21_X1 FSM_U3 ( .B1(FSM_n87), .B2(FSM_n88), .A(FSM_n29), .ZN(FSM_n82) );
  DFF_X1 FSM_LFSR_reg_5_ ( .D(FSM_n71), .CK(CLK), .Q(FSM_n27), .QN(FSM_n10) );
  DFF_X1 FSM_CONST_reg_0_ ( .D(FSM_CONST_internal[0]), .CK(CLK), .Q(CONST[0]), 
        .QN() );
  DFF_X1 FSM_CONST_reg_3_ ( .D(FSM_CONST_internal_3), .CK(CLK), .Q(CONST[3]), 
        .QN() );
  DFF_X1 FSM_CONST_reg_1_ ( .D(FSM_CONST_internal[1]), .CK(CLK), .Q(CONST[1]), 
        .QN() );
  DFF_X1 FSM_CONST_reg_7_ ( .D(FSM_CONST_internal_7), .CK(CLK), .Q(CONST[7]), 
        .QN() );
  DFF_X1 FSM_STATE_reg_1_ ( .D(FSM_n78), .CK(CLK), .Q(), .QN(FSM_n17) );
  DFF_X1 FSM_LFSR_reg_6_ ( .D(FSM_n70), .CK(CLK), .Q(FSM_n23), .QN(FSM_n8) );
  DFF_X1 FSM_LFSR_reg_4_ ( .D(FSM_n72), .CK(CLK), .Q(FSM_n22), .QN(FSM_n11) );
  DFF_X1 FSM_LFSR_reg_3_ ( .D(FSM_n73), .CK(CLK), .Q(FSM_n20), .QN(FSM_n12) );
  DFF_X1 FSM_LFSR_reg_2_ ( .D(FSM_n74), .CK(CLK), .Q(FSM_n21), .QN(FSM_n13) );
  DFF_X1 FSM_LFSR_reg_1_ ( .D(FSM_n75), .CK(CLK), .Q(FSM_n24), .QN(FSM_n14) );
  DFF_X1 FSM_LFSR_reg_0_ ( .D(FSM_n76), .CK(CLK), .Q(FSM_n25), .QN(FSM_n15) );
  DFF_X1 FSM_LFSR_reg_7_ ( .D(FSM_n77), .CK(CLK), .Q(FSM_n26), .QN(FSM_n7) );
  DFF_X1 FSM_STATE_reg_2_ ( .D(FSM_n1), .CK(CLK), .Q(FSM_n87), .QN() );
  DFF_X1 FSM_STATE_reg_0_ ( .D(FSM_n79), .CK(CLK), .Q(FSM_n28), .QN(FSM_n18)
         );
endmodule

