
module circuit ( clk, reset, input_s1, input_s2, input_s3, r, output_s1, 
        output_s2, output_s3, Key1, Key2, Key3, enc_dec, done );
  input [63:0] input_s1;
  input [63:0] input_s2;
  input [63:0] input_s3;
  input [69:0] r;
  output [63:0] output_s1;
  output [63:0] output_s2;
  output [63:0] output_s3;
  input [127:0] Key1;
  input [127:0] Key2;
  input [127:0] Key3;
  input clk, reset, enc_dec;
  output done;
  wire   roundHalf_Select_Signal, roundEnd_Select_Signal, MyController_n36,
         MyController_n35, MyController_n34, MyController_n33,
         MyController_n32, MyController_n31, MyController_n29,
         MyController_n28, MyController_n27, MyController_n26,
         MyController_n25, MyController_n24, MyController_n23,
         MyController_n22, MyController_n21, MyController_n20,
         MyController_n19, MyController_n18, MyController_n17,
         MyController_n16, MyController_n15, MyController_n14,
         MyController_n13, MyController_n12, MyController_n11,
         MyController_n10, MyController_n9, MyController_n8, MyController_n7,
         MyController_n6, MyController_n5, MyController_n3, MyController_n2,
         MyController_n47, MyController_n46, MyController_n45,
         MyController_n44, MyController_n43, MyController_n4, MyController_n77,
         MyController_n76, MyController_n75, MyController_n74,
         MyController_n40, MyController_n38, MyController_n30,
         MyController_N27, MyController_N25, MyController_N19,
         MyController_N18, MyController_N17, prince_n3,
         prince_selected_Key3_0_, prince_selected_Key3_1_,
         prince_selected_Key3_2_, prince_selected_Key3_3_,
         prince_selected_Key3_4_, prince_selected_Key3_5_,
         prince_selected_Key3_6_, prince_selected_Key3_7_,
         prince_selected_Key3_8_, prince_selected_Key3_9_,
         prince_selected_Key3_10_, prince_selected_Key3_11_,
         prince_selected_Key3_12_, prince_selected_Key3_13_,
         prince_selected_Key3_14_, prince_selected_Key3_15_,
         prince_selected_Key3_16_, prince_selected_Key3_17_,
         prince_selected_Key3_18_, prince_selected_Key3_19_,
         prince_selected_Key3_20_, prince_selected_Key3_21_,
         prince_selected_Key3_22_, prince_selected_Key3_23_,
         prince_selected_Key3_24_, prince_selected_Key3_25_,
         prince_selected_Key3_26_, prince_selected_Key3_27_,
         prince_selected_Key3_28_, prince_selected_Key3_29_,
         prince_selected_Key3_30_, prince_selected_Key3_31_,
         prince_selected_Key3_32_, prince_selected_Key3_33_,
         prince_selected_Key3_34_, prince_selected_Key3_35_,
         prince_selected_Key3_36_, prince_selected_Key3_37_,
         prince_selected_Key3_38_, prince_selected_Key3_39_,
         prince_selected_Key3_40_, prince_selected_Key3_41_,
         prince_selected_Key3_42_, prince_selected_Key3_43_,
         prince_selected_Key3_44_, prince_selected_Key3_45_,
         prince_selected_Key3_46_, prince_selected_Key3_47_,
         prince_selected_Key3_48_, prince_selected_Key3_49_,
         prince_selected_Key3_50_, prince_selected_Key3_51_,
         prince_selected_Key3_52_, prince_selected_Key3_53_,
         prince_selected_Key3_54_, prince_selected_Key3_55_,
         prince_selected_Key3_56_, prince_selected_Key3_57_,
         prince_selected_Key3_58_, prince_selected_Key3_59_,
         prince_selected_Key3_60_, prince_selected_Key3_61_,
         prince_selected_Key3_62_, prince_selected_Key3_63_,
         prince_selected_Key2_0_, prince_selected_Key2_1_,
         prince_selected_Key2_2_, prince_selected_Key2_3_,
         prince_selected_Key2_4_, prince_selected_Key2_5_,
         prince_selected_Key2_6_, prince_selected_Key2_7_,
         prince_selected_Key2_8_, prince_selected_Key2_9_,
         prince_selected_Key2_10_, prince_selected_Key2_11_,
         prince_selected_Key2_12_, prince_selected_Key2_13_,
         prince_selected_Key2_14_, prince_selected_Key2_15_,
         prince_selected_Key2_16_, prince_selected_Key2_17_,
         prince_selected_Key2_18_, prince_selected_Key2_19_,
         prince_selected_Key2_20_, prince_selected_Key2_21_,
         prince_selected_Key2_22_, prince_selected_Key2_23_,
         prince_selected_Key2_24_, prince_selected_Key2_25_,
         prince_selected_Key2_26_, prince_selected_Key2_27_,
         prince_selected_Key2_28_, prince_selected_Key2_29_,
         prince_selected_Key2_30_, prince_selected_Key2_31_,
         prince_selected_Key2_32_, prince_selected_Key2_33_,
         prince_selected_Key2_34_, prince_selected_Key2_35_,
         prince_selected_Key2_36_, prince_selected_Key2_37_,
         prince_selected_Key2_38_, prince_selected_Key2_39_,
         prince_selected_Key2_40_, prince_selected_Key2_41_,
         prince_selected_Key2_42_, prince_selected_Key2_43_,
         prince_selected_Key2_44_, prince_selected_Key2_45_,
         prince_selected_Key2_46_, prince_selected_Key2_47_,
         prince_selected_Key2_48_, prince_selected_Key2_49_,
         prince_selected_Key2_50_, prince_selected_Key2_51_,
         prince_selected_Key2_52_, prince_selected_Key2_53_,
         prince_selected_Key2_54_, prince_selected_Key2_55_,
         prince_selected_Key2_56_, prince_selected_Key2_57_,
         prince_selected_Key2_58_, prince_selected_Key2_59_,
         prince_selected_Key2_60_, prince_selected_Key2_61_,
         prince_selected_Key2_62_, prince_selected_Key2_63_,
         prince_selected_Key1_0_, prince_selected_Key1_1_,
         prince_selected_Key1_2_, prince_selected_Key1_3_,
         prince_selected_Key1_4_, prince_selected_Key1_5_,
         prince_selected_Key1_6_, prince_selected_Key1_7_,
         prince_selected_Key1_8_, prince_selected_Key1_9_,
         prince_selected_Key1_10_, prince_selected_Key1_11_,
         prince_selected_Key1_12_, prince_selected_Key1_13_,
         prince_selected_Key1_14_, prince_selected_Key1_15_,
         prince_selected_Key1_16_, prince_selected_Key1_17_,
         prince_selected_Key1_18_, prince_selected_Key1_19_,
         prince_selected_Key1_20_, prince_selected_Key1_21_,
         prince_selected_Key1_22_, prince_selected_Key1_23_,
         prince_selected_Key1_24_, prince_selected_Key1_25_,
         prince_selected_Key1_26_, prince_selected_Key1_27_,
         prince_selected_Key1_28_, prince_selected_Key1_29_,
         prince_selected_Key1_30_, prince_selected_Key1_31_,
         prince_selected_Key1_32_, prince_selected_Key1_33_,
         prince_selected_Key1_34_, prince_selected_Key1_35_,
         prince_selected_Key1_36_, prince_selected_Key1_37_,
         prince_selected_Key1_38_, prince_selected_Key1_39_,
         prince_selected_Key1_40_, prince_selected_Key1_41_,
         prince_selected_Key1_42_, prince_selected_Key1_43_,
         prince_selected_Key1_44_, prince_selected_Key1_45_,
         prince_selected_Key1_46_, prince_selected_Key1_47_,
         prince_selected_Key1_48_, prince_selected_Key1_49_,
         prince_selected_Key1_50_, prince_selected_Key1_51_,
         prince_selected_Key1_52_, prince_selected_Key1_53_,
         prince_selected_Key1_54_, prince_selected_Key1_55_,
         prince_selected_Key1_56_, prince_selected_Key1_57_,
         prince_selected_Key1_58_, prince_selected_Key1_59_,
         prince_selected_Key1_60_, prince_selected_Key1_61_,
         prince_selected_Key1_62_, prince_selected_Key1_63_,
         prince_enc_dec_xor_reset, prince_k_0_p_share3_0_,
         prince_k_0_p_share2_0_, prince_k_0_p_share1_0_, prince_KeyMUX1_n10,
         prince_KeyMUX1_n9, prince_KeyMUX1_n8, prince_KeyMUX1_n7,
         prince_KeyMUX2_n10, prince_KeyMUX2_n9, prince_KeyMUX2_n8,
         prince_KeyMUX2_n7, prince_KeyMUX3_n9, prince_KeyMUX3_n8,
         prince_KeyMUX3_n7, prince_AddKey1_XORInst_0_0_n3,
         prince_AddKey1_XORInst_0_1_n3, prince_AddKey1_XORInst_0_2_n3,
         prince_AddKey1_XORInst_0_3_n3, prince_AddKey1_XORInst_1_0_n3,
         prince_AddKey1_XORInst_1_1_n3, prince_AddKey1_XORInst_1_2_n3,
         prince_AddKey1_XORInst_1_3_n3, prince_AddKey1_XORInst_2_0_n3,
         prince_AddKey1_XORInst_2_1_n3, prince_AddKey1_XORInst_2_2_n3,
         prince_AddKey1_XORInst_2_3_n3, prince_AddKey1_XORInst_3_0_n3,
         prince_AddKey1_XORInst_3_1_n3, prince_AddKey1_XORInst_3_2_n3,
         prince_AddKey1_XORInst_3_3_n3, prince_AddKey1_XORInst_4_0_n3,
         prince_AddKey1_XORInst_4_1_n3, prince_AddKey1_XORInst_4_2_n3,
         prince_AddKey1_XORInst_4_3_n3, prince_AddKey1_XORInst_5_0_n3,
         prince_AddKey1_XORInst_5_1_n3, prince_AddKey1_XORInst_5_2_n3,
         prince_AddKey1_XORInst_5_3_n3, prince_AddKey1_XORInst_6_0_n3,
         prince_AddKey1_XORInst_6_1_n3, prince_AddKey1_XORInst_6_2_n3,
         prince_AddKey1_XORInst_6_3_n3, prince_AddKey1_XORInst_7_0_n3,
         prince_AddKey1_XORInst_7_1_n3, prince_AddKey1_XORInst_7_2_n3,
         prince_AddKey1_XORInst_7_3_n3, prince_AddKey1_XORInst_8_0_n3,
         prince_AddKey1_XORInst_8_1_n3, prince_AddKey1_XORInst_8_2_n3,
         prince_AddKey1_XORInst_8_3_n3, prince_AddKey1_XORInst_9_0_n3,
         prince_AddKey1_XORInst_9_1_n3, prince_AddKey1_XORInst_9_2_n3,
         prince_AddKey1_XORInst_9_3_n3, prince_AddKey1_XORInst_10_0_n3,
         prince_AddKey1_XORInst_10_1_n3, prince_AddKey1_XORInst_10_2_n3,
         prince_AddKey1_XORInst_10_3_n3, prince_AddKey1_XORInst_11_0_n3,
         prince_AddKey1_XORInst_11_1_n3, prince_AddKey1_XORInst_11_2_n3,
         prince_AddKey1_XORInst_11_3_n3, prince_AddKey1_XORInst_12_0_n3,
         prince_AddKey1_XORInst_12_1_n3, prince_AddKey1_XORInst_12_2_n3,
         prince_AddKey1_XORInst_12_3_n3, prince_AddKey1_XORInst_13_0_n3,
         prince_AddKey1_XORInst_13_1_n3, prince_AddKey1_XORInst_13_2_n3,
         prince_AddKey1_XORInst_13_3_n3, prince_AddKey1_XORInst_14_0_n3,
         prince_AddKey1_XORInst_14_1_n3, prince_AddKey1_XORInst_14_2_n3,
         prince_AddKey1_XORInst_14_3_n3, prince_AddKey1_XORInst_15_0_n3,
         prince_AddKey1_XORInst_15_1_n3, prince_AddKey1_XORInst_15_2_n3,
         prince_AddKey1_XORInst_15_3_n3, prince_AddKey2_XORInst_0_0_n3,
         prince_AddKey2_XORInst_0_1_n3, prince_AddKey2_XORInst_0_2_n3,
         prince_AddKey2_XORInst_0_3_n3, prince_AddKey2_XORInst_1_0_n3,
         prince_AddKey2_XORInst_1_1_n3, prince_AddKey2_XORInst_1_2_n3,
         prince_AddKey2_XORInst_1_3_n3, prince_AddKey2_XORInst_2_0_n3,
         prince_AddKey2_XORInst_2_1_n3, prince_AddKey2_XORInst_2_2_n3,
         prince_AddKey2_XORInst_2_3_n3, prince_AddKey2_XORInst_3_0_n3,
         prince_AddKey2_XORInst_3_1_n3, prince_AddKey2_XORInst_3_2_n3,
         prince_AddKey2_XORInst_3_3_n3, prince_AddKey2_XORInst_4_0_n3,
         prince_AddKey2_XORInst_4_1_n3, prince_AddKey2_XORInst_4_2_n3,
         prince_AddKey2_XORInst_4_3_n3, prince_AddKey2_XORInst_5_0_n3,
         prince_AddKey2_XORInst_5_1_n3, prince_AddKey2_XORInst_5_2_n3,
         prince_AddKey2_XORInst_5_3_n3, prince_AddKey2_XORInst_6_0_n3,
         prince_AddKey2_XORInst_6_1_n3, prince_AddKey2_XORInst_6_2_n3,
         prince_AddKey2_XORInst_6_3_n3, prince_AddKey2_XORInst_7_0_n3,
         prince_AddKey2_XORInst_7_1_n3, prince_AddKey2_XORInst_7_2_n3,
         prince_AddKey2_XORInst_7_3_n3, prince_AddKey2_XORInst_8_0_n3,
         prince_AddKey2_XORInst_8_1_n3, prince_AddKey2_XORInst_8_2_n3,
         prince_AddKey2_XORInst_8_3_n3, prince_AddKey2_XORInst_9_0_n3,
         prince_AddKey2_XORInst_9_1_n3, prince_AddKey2_XORInst_9_2_n3,
         prince_AddKey2_XORInst_9_3_n3, prince_AddKey2_XORInst_10_0_n3,
         prince_AddKey2_XORInst_10_1_n3, prince_AddKey2_XORInst_10_2_n3,
         prince_AddKey2_XORInst_10_3_n3, prince_AddKey2_XORInst_11_0_n3,
         prince_AddKey2_XORInst_11_1_n3, prince_AddKey2_XORInst_11_2_n3,
         prince_AddKey2_XORInst_11_3_n3, prince_AddKey2_XORInst_12_0_n3,
         prince_AddKey2_XORInst_12_1_n3, prince_AddKey2_XORInst_12_2_n3,
         prince_AddKey2_XORInst_12_3_n3, prince_AddKey2_XORInst_13_0_n3,
         prince_AddKey2_XORInst_13_1_n3, prince_AddKey2_XORInst_13_2_n3,
         prince_AddKey2_XORInst_13_3_n3, prince_AddKey2_XORInst_14_0_n3,
         prince_AddKey2_XORInst_14_1_n3, prince_AddKey2_XORInst_14_2_n3,
         prince_AddKey2_XORInst_14_3_n3, prince_AddKey2_XORInst_15_0_n3,
         prince_AddKey2_XORInst_15_1_n3, prince_AddKey2_XORInst_15_2_n3,
         prince_AddKey2_XORInst_15_3_n3, prince_AddKey3_XORInst_0_0_n3,
         prince_AddKey3_XORInst_0_1_n3, prince_AddKey3_XORInst_0_2_n3,
         prince_AddKey3_XORInst_0_3_n3, prince_AddKey3_XORInst_1_0_n3,
         prince_AddKey3_XORInst_1_1_n3, prince_AddKey3_XORInst_1_2_n3,
         prince_AddKey3_XORInst_1_3_n3, prince_AddKey3_XORInst_2_0_n3,
         prince_AddKey3_XORInst_2_1_n3, prince_AddKey3_XORInst_2_2_n3,
         prince_AddKey3_XORInst_2_3_n3, prince_AddKey3_XORInst_3_0_n3,
         prince_AddKey3_XORInst_3_1_n3, prince_AddKey3_XORInst_3_2_n3,
         prince_AddKey3_XORInst_3_3_n3, prince_AddKey3_XORInst_4_0_n3,
         prince_AddKey3_XORInst_4_1_n3, prince_AddKey3_XORInst_4_2_n3,
         prince_AddKey3_XORInst_4_3_n3, prince_AddKey3_XORInst_5_0_n3,
         prince_AddKey3_XORInst_5_1_n3, prince_AddKey3_XORInst_5_2_n3,
         prince_AddKey3_XORInst_5_3_n3, prince_AddKey3_XORInst_6_0_n3,
         prince_AddKey3_XORInst_6_1_n3, prince_AddKey3_XORInst_6_2_n3,
         prince_AddKey3_XORInst_6_3_n3, prince_AddKey3_XORInst_7_0_n3,
         prince_AddKey3_XORInst_7_1_n3, prince_AddKey3_XORInst_7_2_n3,
         prince_AddKey3_XORInst_7_3_n3, prince_AddKey3_XORInst_8_0_n3,
         prince_AddKey3_XORInst_8_1_n3, prince_AddKey3_XORInst_8_2_n3,
         prince_AddKey3_XORInst_8_3_n3, prince_AddKey3_XORInst_9_0_n3,
         prince_AddKey3_XORInst_9_1_n3, prince_AddKey3_XORInst_9_2_n3,
         prince_AddKey3_XORInst_9_3_n3, prince_AddKey3_XORInst_10_0_n3,
         prince_AddKey3_XORInst_10_1_n3, prince_AddKey3_XORInst_10_2_n3,
         prince_AddKey3_XORInst_10_3_n3, prince_AddKey3_XORInst_11_0_n3,
         prince_AddKey3_XORInst_11_1_n3, prince_AddKey3_XORInst_11_2_n3,
         prince_AddKey3_XORInst_11_3_n3, prince_AddKey3_XORInst_12_0_n3,
         prince_AddKey3_XORInst_12_1_n3, prince_AddKey3_XORInst_12_2_n3,
         prince_AddKey3_XORInst_12_3_n3, prince_AddKey3_XORInst_13_0_n3,
         prince_AddKey3_XORInst_13_1_n3, prince_AddKey3_XORInst_13_2_n3,
         prince_AddKey3_XORInst_13_3_n3, prince_AddKey3_XORInst_14_0_n3,
         prince_AddKey3_XORInst_14_1_n3, prince_AddKey3_XORInst_14_2_n3,
         prince_AddKey3_XORInst_14_3_n3, prince_AddKey3_XORInst_15_0_n3,
         prince_AddKey3_XORInst_15_1_n3, prince_AddKey3_XORInst_15_2_n3,
         prince_AddKey3_XORInst_15_3_n3, prince_rounds_n65, prince_rounds_n64,
         prince_rounds_n63, prince_rounds_n62, prince_rounds_n61,
         prince_rounds_n60, prince_rounds_n59, prince_rounds_n58,
         prince_rounds_n57, prince_rounds_n56, prince_rounds_n55,
         prince_rounds_n54, prince_rounds_n53, prince_rounds_n52,
         prince_rounds_n51, prince_rounds_n50, prince_rounds_n49,
         prince_rounds_n48, prince_rounds_n47, prince_rounds_n46,
         prince_rounds_n45, prince_rounds_n44, prince_rounds_n43,
         prince_rounds_n42, prince_rounds_n41, prince_rounds_n40,
         prince_rounds_n39, prince_rounds_n38, prince_rounds_n37,
         prince_rounds_n36, prince_rounds_n35, prince_rounds_n34,
         prince_rounds_n33, prince_rounds_n32, prince_rounds_n31,
         prince_rounds_n30, prince_rounds_n29, prince_rounds_n28,
         prince_rounds_n27, prince_rounds_n26, prince_rounds_n25,
         prince_rounds_n24, prince_rounds_n23, prince_rounds_n22,
         prince_rounds_n21, prince_rounds_n20, prince_rounds_n19,
         prince_rounds_n18, prince_rounds_k1_XOR_round_Constant_0_,
         prince_rounds_k1_XOR_round_Constant_1_,
         prince_rounds_k1_XOR_round_Constant_2_,
         prince_rounds_k1_XOR_round_Constant_3_,
         prince_rounds_k1_XOR_round_Constant_4_,
         prince_rounds_k1_XOR_round_Constant_5_,
         prince_rounds_k1_XOR_round_Constant_6_,
         prince_rounds_k1_XOR_round_Constant_7_,
         prince_rounds_k1_XOR_round_Constant_8_,
         prince_rounds_k1_XOR_round_Constant_9_,
         prince_rounds_k1_XOR_round_Constant_10_,
         prince_rounds_k1_XOR_round_Constant_11_,
         prince_rounds_k1_XOR_round_Constant_12_,
         prince_rounds_k1_XOR_round_Constant_13_,
         prince_rounds_k1_XOR_round_Constant_14_,
         prince_rounds_k1_XOR_round_Constant_15_,
         prince_rounds_k1_XOR_round_Constant_16_,
         prince_rounds_k1_XOR_round_Constant_17_,
         prince_rounds_k1_XOR_round_Constant_18_,
         prince_rounds_k1_XOR_round_Constant_19_,
         prince_rounds_k1_XOR_round_Constant_20_,
         prince_rounds_k1_XOR_round_Constant_21_,
         prince_rounds_k1_XOR_round_Constant_22_,
         prince_rounds_k1_XOR_round_Constant_23_,
         prince_rounds_k1_XOR_round_Constant_24_,
         prince_rounds_k1_XOR_round_Constant_25_,
         prince_rounds_k1_XOR_round_Constant_26_,
         prince_rounds_k1_XOR_round_Constant_27_,
         prince_rounds_k1_XOR_round_Constant_28_,
         prince_rounds_k1_XOR_round_Constant_29_,
         prince_rounds_k1_XOR_round_Constant_30_,
         prince_rounds_k1_XOR_round_Constant_31_,
         prince_rounds_k1_XOR_round_Constant_32_,
         prince_rounds_k1_XOR_round_Constant_33_,
         prince_rounds_k1_XOR_round_Constant_34_,
         prince_rounds_k1_XOR_round_Constant_35_,
         prince_rounds_k1_XOR_round_Constant_36_,
         prince_rounds_k1_XOR_round_Constant_37_,
         prince_rounds_k1_XOR_round_Constant_38_,
         prince_rounds_k1_XOR_round_Constant_39_,
         prince_rounds_k1_XOR_round_Constant_40_,
         prince_rounds_k1_XOR_round_Constant_41_,
         prince_rounds_k1_XOR_round_Constant_42_,
         prince_rounds_k1_XOR_round_Constant_43_,
         prince_rounds_k1_XOR_round_Constant_44_,
         prince_rounds_k1_XOR_round_Constant_45_,
         prince_rounds_k1_XOR_round_Constant_46_,
         prince_rounds_k1_XOR_round_Constant_47_,
         prince_rounds_k1_XOR_round_Constant_48_,
         prince_rounds_k1_XOR_round_Constant_49_,
         prince_rounds_k1_XOR_round_Constant_50_,
         prince_rounds_k1_XOR_round_Constant_51_,
         prince_rounds_k1_XOR_round_Constant_52_,
         prince_rounds_k1_XOR_round_Constant_53_,
         prince_rounds_k1_XOR_round_Constant_54_,
         prince_rounds_k1_XOR_round_Constant_55_,
         prince_rounds_k1_XOR_round_Constant_56_,
         prince_rounds_k1_XOR_round_Constant_57_,
         prince_rounds_k1_XOR_round_Constant_58_,
         prince_rounds_k1_XOR_round_Constant_59_,
         prince_rounds_k1_XOR_round_Constant_60_,
         prince_rounds_k1_XOR_round_Constant_61_,
         prince_rounds_k1_XOR_round_Constant_62_,
         prince_rounds_k1_XOR_round_Constant_63_,
         prince_rounds_constant_MUX_n46, prince_rounds_constant_MUX_n45,
         prince_rounds_constant_MUX_n44, prince_rounds_constant_MUX_n43,
         prince_rounds_constant_MUX_n42, prince_rounds_constant_MUX_n41,
         prince_rounds_constant_MUX_n40, prince_rounds_constant_MUX_n39,
         prince_rounds_constant_MUX_n38, prince_rounds_constant_MUX_n37,
         prince_rounds_constant_MUX_n36, prince_rounds_constant_MUX_n35,
         prince_rounds_constant_MUX_n34, prince_rounds_constant_MUX_n33,
         prince_rounds_constant_MUX_n32, prince_rounds_constant_MUX_n31,
         prince_rounds_constant_MUX_n30, prince_rounds_constant_MUX_n29,
         prince_rounds_constant_MUX_n28, prince_rounds_constant_MUX_n27,
         prince_rounds_constant_MUX_n26, prince_rounds_constant_MUX_n25,
         prince_rounds_constant_MUX_n24, prince_rounds_constant_MUX_n23,
         prince_rounds_constant_MUX_n22, prince_rounds_constant_MUX_n21,
         prince_rounds_constant_MUX_n20, prince_rounds_constant_MUX_n19,
         prince_rounds_constant_MUX_n18, prince_rounds_constant_MUX_n17,
         prince_rounds_constant_MUX_n16, prince_rounds_constant_MUX_n15,
         prince_rounds_constant_MUX_n14, prince_rounds_constant_MUX_n13,
         prince_rounds_constant_MUX_n12, prince_rounds_constant_MUX_n11,
         prince_rounds_constant_MUX_n10, prince_rounds_constant_MUX_n9,
         prince_rounds_constant_MUX_n8, prince_rounds_constant_MUX_n7,
         prince_rounds_constant_MUX_n6, prince_rounds_constant_MUX_n5,
         prince_rounds_constant_MUX_n4, prince_rounds_constant_MUX_n3,
         prince_rounds_constant_MUX_n2, prince_rounds_constant_MUX_n1,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_0_0_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_0_1_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_0_2_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_0_3_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_1_0_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_1_1_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_1_2_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_1_3_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_2_0_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_2_1_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_2_2_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_2_3_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_3_0_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_3_1_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_3_2_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_3_3_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_4_0_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_4_1_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_4_2_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_4_3_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_5_0_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_5_1_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_5_2_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_5_3_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_6_0_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_6_1_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_6_2_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_6_3_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_7_0_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_7_1_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_7_2_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_7_3_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_8_0_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_8_1_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_8_2_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_8_3_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_9_0_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_9_1_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_9_2_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_9_3_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_10_0_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_10_1_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_10_2_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_10_3_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_11_0_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_11_1_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_11_2_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_11_3_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_12_0_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_12_1_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_12_2_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_12_3_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_13_0_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_13_1_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_13_2_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_13_3_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_14_0_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_14_1_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_14_2_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_14_3_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_15_0_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_15_1_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_15_2_n3,
         prince_rounds_k1_XOR_round_Constant_module_XORInst_15_3_n3,
         prince_rounds_AddKey1_XORInst_0_0_n3,
         prince_rounds_AddKey1_XORInst_0_1_n3,
         prince_rounds_AddKey1_XORInst_0_2_n3,
         prince_rounds_AddKey1_XORInst_0_3_n3,
         prince_rounds_AddKey1_XORInst_1_0_n3,
         prince_rounds_AddKey1_XORInst_1_1_n3,
         prince_rounds_AddKey1_XORInst_1_2_n3,
         prince_rounds_AddKey1_XORInst_1_3_n3,
         prince_rounds_AddKey1_XORInst_2_0_n3,
         prince_rounds_AddKey1_XORInst_2_1_n3,
         prince_rounds_AddKey1_XORInst_2_2_n3,
         prince_rounds_AddKey1_XORInst_2_3_n3,
         prince_rounds_AddKey1_XORInst_3_0_n3,
         prince_rounds_AddKey1_XORInst_3_1_n3,
         prince_rounds_AddKey1_XORInst_3_2_n3,
         prince_rounds_AddKey1_XORInst_3_3_n3,
         prince_rounds_AddKey1_XORInst_4_0_n3,
         prince_rounds_AddKey1_XORInst_4_1_n3,
         prince_rounds_AddKey1_XORInst_4_2_n3,
         prince_rounds_AddKey1_XORInst_4_3_n3,
         prince_rounds_AddKey1_XORInst_5_0_n3,
         prince_rounds_AddKey1_XORInst_5_1_n3,
         prince_rounds_AddKey1_XORInst_5_2_n3,
         prince_rounds_AddKey1_XORInst_5_3_n3,
         prince_rounds_AddKey1_XORInst_6_0_n3,
         prince_rounds_AddKey1_XORInst_6_1_n3,
         prince_rounds_AddKey1_XORInst_6_2_n3,
         prince_rounds_AddKey1_XORInst_6_3_n3,
         prince_rounds_AddKey1_XORInst_7_0_n3,
         prince_rounds_AddKey1_XORInst_7_1_n3,
         prince_rounds_AddKey1_XORInst_7_2_n3,
         prince_rounds_AddKey1_XORInst_7_3_n3,
         prince_rounds_AddKey1_XORInst_8_0_n3,
         prince_rounds_AddKey1_XORInst_8_1_n3,
         prince_rounds_AddKey1_XORInst_8_2_n3,
         prince_rounds_AddKey1_XORInst_8_3_n3,
         prince_rounds_AddKey1_XORInst_9_0_n3,
         prince_rounds_AddKey1_XORInst_9_1_n3,
         prince_rounds_AddKey1_XORInst_9_2_n3,
         prince_rounds_AddKey1_XORInst_9_3_n3,
         prince_rounds_AddKey1_XORInst_10_0_n3,
         prince_rounds_AddKey1_XORInst_10_1_n3,
         prince_rounds_AddKey1_XORInst_10_2_n3,
         prince_rounds_AddKey1_XORInst_10_3_n3,
         prince_rounds_AddKey1_XORInst_11_0_n3,
         prince_rounds_AddKey1_XORInst_11_1_n3,
         prince_rounds_AddKey1_XORInst_11_2_n3,
         prince_rounds_AddKey1_XORInst_11_3_n3,
         prince_rounds_AddKey1_XORInst_12_0_n3,
         prince_rounds_AddKey1_XORInst_12_1_n3,
         prince_rounds_AddKey1_XORInst_12_2_n3,
         prince_rounds_AddKey1_XORInst_12_3_n3,
         prince_rounds_AddKey1_XORInst_13_0_n3,
         prince_rounds_AddKey1_XORInst_13_1_n3,
         prince_rounds_AddKey1_XORInst_13_2_n3,
         prince_rounds_AddKey1_XORInst_13_3_n3,
         prince_rounds_AddKey1_XORInst_14_0_n3,
         prince_rounds_AddKey1_XORInst_14_1_n3,
         prince_rounds_AddKey1_XORInst_14_2_n3,
         prince_rounds_AddKey1_XORInst_14_3_n3,
         prince_rounds_AddKey1_XORInst_15_0_n3,
         prince_rounds_AddKey1_XORInst_15_1_n3,
         prince_rounds_AddKey1_XORInst_15_2_n3,
         prince_rounds_AddKey1_XORInst_15_3_n3,
         prince_rounds_AddKey2_XORInst_0_0_n3,
         prince_rounds_AddKey2_XORInst_0_1_n3,
         prince_rounds_AddKey2_XORInst_0_2_n3,
         prince_rounds_AddKey2_XORInst_0_3_n3,
         prince_rounds_AddKey2_XORInst_1_0_n3,
         prince_rounds_AddKey2_XORInst_1_1_n3,
         prince_rounds_AddKey2_XORInst_1_2_n3,
         prince_rounds_AddKey2_XORInst_1_3_n3,
         prince_rounds_AddKey2_XORInst_2_0_n3,
         prince_rounds_AddKey2_XORInst_2_1_n3,
         prince_rounds_AddKey2_XORInst_2_2_n3,
         prince_rounds_AddKey2_XORInst_2_3_n3,
         prince_rounds_AddKey2_XORInst_3_0_n3,
         prince_rounds_AddKey2_XORInst_3_1_n3,
         prince_rounds_AddKey2_XORInst_3_2_n3,
         prince_rounds_AddKey2_XORInst_3_3_n3,
         prince_rounds_AddKey2_XORInst_4_0_n3,
         prince_rounds_AddKey2_XORInst_4_1_n3,
         prince_rounds_AddKey2_XORInst_4_2_n3,
         prince_rounds_AddKey2_XORInst_4_3_n3,
         prince_rounds_AddKey2_XORInst_5_0_n3,
         prince_rounds_AddKey2_XORInst_5_1_n3,
         prince_rounds_AddKey2_XORInst_5_2_n3,
         prince_rounds_AddKey2_XORInst_5_3_n3,
         prince_rounds_AddKey2_XORInst_6_0_n3,
         prince_rounds_AddKey2_XORInst_6_1_n3,
         prince_rounds_AddKey2_XORInst_6_2_n3,
         prince_rounds_AddKey2_XORInst_6_3_n3,
         prince_rounds_AddKey2_XORInst_7_0_n3,
         prince_rounds_AddKey2_XORInst_7_1_n3,
         prince_rounds_AddKey2_XORInst_7_2_n3,
         prince_rounds_AddKey2_XORInst_7_3_n3,
         prince_rounds_AddKey2_XORInst_8_0_n3,
         prince_rounds_AddKey2_XORInst_8_1_n3,
         prince_rounds_AddKey2_XORInst_8_2_n3,
         prince_rounds_AddKey2_XORInst_8_3_n3,
         prince_rounds_AddKey2_XORInst_9_0_n3,
         prince_rounds_AddKey2_XORInst_9_1_n3,
         prince_rounds_AddKey2_XORInst_9_2_n3,
         prince_rounds_AddKey2_XORInst_9_3_n3,
         prince_rounds_AddKey2_XORInst_10_0_n3,
         prince_rounds_AddKey2_XORInst_10_1_n3,
         prince_rounds_AddKey2_XORInst_10_2_n3,
         prince_rounds_AddKey2_XORInst_10_3_n3,
         prince_rounds_AddKey2_XORInst_11_0_n3,
         prince_rounds_AddKey2_XORInst_11_1_n3,
         prince_rounds_AddKey2_XORInst_11_2_n3,
         prince_rounds_AddKey2_XORInst_11_3_n3,
         prince_rounds_AddKey2_XORInst_12_0_n3,
         prince_rounds_AddKey2_XORInst_12_1_n3,
         prince_rounds_AddKey2_XORInst_12_2_n3,
         prince_rounds_AddKey2_XORInst_12_3_n3,
         prince_rounds_AddKey2_XORInst_13_0_n3,
         prince_rounds_AddKey2_XORInst_13_1_n3,
         prince_rounds_AddKey2_XORInst_13_2_n3,
         prince_rounds_AddKey2_XORInst_13_3_n3,
         prince_rounds_AddKey2_XORInst_14_0_n3,
         prince_rounds_AddKey2_XORInst_14_1_n3,
         prince_rounds_AddKey2_XORInst_14_2_n3,
         prince_rounds_AddKey2_XORInst_14_3_n3,
         prince_rounds_AddKey2_XORInst_15_0_n3,
         prince_rounds_AddKey2_XORInst_15_1_n3,
         prince_rounds_AddKey2_XORInst_15_2_n3,
         prince_rounds_AddKey2_XORInst_15_3_n3,
         prince_rounds_AddKey3_XORInst_0_0_n3,
         prince_rounds_AddKey3_XORInst_0_1_n3,
         prince_rounds_AddKey3_XORInst_0_2_n3,
         prince_rounds_AddKey3_XORInst_0_3_n3,
         prince_rounds_AddKey3_XORInst_1_0_n3,
         prince_rounds_AddKey3_XORInst_1_1_n3,
         prince_rounds_AddKey3_XORInst_1_2_n3,
         prince_rounds_AddKey3_XORInst_1_3_n3,
         prince_rounds_AddKey3_XORInst_2_0_n3,
         prince_rounds_AddKey3_XORInst_2_1_n3,
         prince_rounds_AddKey3_XORInst_2_2_n3,
         prince_rounds_AddKey3_XORInst_2_3_n3,
         prince_rounds_AddKey3_XORInst_3_0_n3,
         prince_rounds_AddKey3_XORInst_3_1_n3,
         prince_rounds_AddKey3_XORInst_3_2_n3,
         prince_rounds_AddKey3_XORInst_3_3_n3,
         prince_rounds_AddKey3_XORInst_4_0_n3,
         prince_rounds_AddKey3_XORInst_4_1_n3,
         prince_rounds_AddKey3_XORInst_4_2_n3,
         prince_rounds_AddKey3_XORInst_4_3_n3,
         prince_rounds_AddKey3_XORInst_5_0_n3,
         prince_rounds_AddKey3_XORInst_5_1_n3,
         prince_rounds_AddKey3_XORInst_5_2_n3,
         prince_rounds_AddKey3_XORInst_5_3_n3,
         prince_rounds_AddKey3_XORInst_6_0_n3,
         prince_rounds_AddKey3_XORInst_6_1_n3,
         prince_rounds_AddKey3_XORInst_6_2_n3,
         prince_rounds_AddKey3_XORInst_6_3_n3,
         prince_rounds_AddKey3_XORInst_7_0_n3,
         prince_rounds_AddKey3_XORInst_7_1_n3,
         prince_rounds_AddKey3_XORInst_7_2_n3,
         prince_rounds_AddKey3_XORInst_7_3_n3,
         prince_rounds_AddKey3_XORInst_8_0_n3,
         prince_rounds_AddKey3_XORInst_8_1_n3,
         prince_rounds_AddKey3_XORInst_8_2_n3,
         prince_rounds_AddKey3_XORInst_8_3_n3,
         prince_rounds_AddKey3_XORInst_9_0_n3,
         prince_rounds_AddKey3_XORInst_9_1_n3,
         prince_rounds_AddKey3_XORInst_9_2_n3,
         prince_rounds_AddKey3_XORInst_9_3_n3,
         prince_rounds_AddKey3_XORInst_10_0_n3,
         prince_rounds_AddKey3_XORInst_10_1_n3,
         prince_rounds_AddKey3_XORInst_10_2_n3,
         prince_rounds_AddKey3_XORInst_10_3_n3,
         prince_rounds_AddKey3_XORInst_11_0_n3,
         prince_rounds_AddKey3_XORInst_11_1_n3,
         prince_rounds_AddKey3_XORInst_11_2_n3,
         prince_rounds_AddKey3_XORInst_11_3_n3,
         prince_rounds_AddKey3_XORInst_12_0_n3,
         prince_rounds_AddKey3_XORInst_12_1_n3,
         prince_rounds_AddKey3_XORInst_12_2_n3,
         prince_rounds_AddKey3_XORInst_12_3_n3,
         prince_rounds_AddKey3_XORInst_13_0_n3,
         prince_rounds_AddKey3_XORInst_13_1_n3,
         prince_rounds_AddKey3_XORInst_13_2_n3,
         prince_rounds_AddKey3_XORInst_13_3_n3,
         prince_rounds_AddKey3_XORInst_14_0_n3,
         prince_rounds_AddKey3_XORInst_14_1_n3,
         prince_rounds_AddKey3_XORInst_14_2_n3,
         prince_rounds_AddKey3_XORInst_14_3_n3,
         prince_rounds_AddKey3_XORInst_15_0_n3,
         prince_rounds_AddKey3_XORInst_15_1_n3,
         prince_rounds_AddKey3_XORInst_15_2_n3,
         prince_rounds_AddKey3_XORInst_15_3_n3, prince_rounds_sub_n4,
         prince_rounds_sub_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_InAffin_s3_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_0_InAffin_s2_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_0_InAffin_s1_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s1_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s1_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s3_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s3_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_n1,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_InAffin_s3_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_1_InAffin_s2_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_1_InAffin_s1_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s1_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s1_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s3_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s3_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_InAffin_s3_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_2_InAffin_s2_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_2_InAffin_s1_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s1_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s1_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s3_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s3_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_InAffin_s3_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_3_InAffin_s2_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_3_InAffin_s1_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s1_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s1_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s3_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s3_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_InAffin_s3_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_4_InAffin_s2_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_4_InAffin_s1_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s1_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s1_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s3_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s3_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_InAffin_s3_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_5_InAffin_s2_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_5_InAffin_s1_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s1_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s1_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s3_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s3_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_InAffin_s3_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_6_InAffin_s2_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_6_InAffin_s1_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s1_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s1_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s3_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s3_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_InAffin_s3_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_7_InAffin_s2_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_7_InAffin_s1_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s1_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s1_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s3_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s3_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_InAffin_s3_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_8_InAffin_s2_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_8_InAffin_s1_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s1_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s1_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s3_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s3_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_InAffin_s3_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_9_InAffin_s2_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_9_InAffin_s1_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s1_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s1_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s3_n19,
         prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s3_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_InAffin_s3_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_10_InAffin_s2_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_10_InAffin_s1_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s1_n19,
         prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s1_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s3_n19,
         prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s3_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_InAffin_s3_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_11_InAffin_s2_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_11_InAffin_s1_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s1_n19,
         prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s1_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s3_n19,
         prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s3_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_InAffin_s3_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_12_InAffin_s2_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_12_InAffin_s1_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s1_n19,
         prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s1_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s3_n19,
         prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s3_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_InAffin_s3_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_13_InAffin_s2_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_13_InAffin_s1_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s1_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s1_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s3_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s3_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_InAffin_s3_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_14_InAffin_s2_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_14_InAffin_s1_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s1_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s1_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s3_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s3_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s3_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_InAffin_s3_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_15_InAffin_s2_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_15_InAffin_s1_3_,
         prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s1_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s1_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_n18,
         prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_n17,
         prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_n16,
         prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_n15,
         prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s3_n21,
         prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s3_n20,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_N1,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_N0,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_0__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_1__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_1__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_2__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_2__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_3__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_4__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_4__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_5__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_5__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_6__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_7__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_7__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_8__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_8__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_9__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_10__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_10__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_11__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_11__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_12__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_13__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_13__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_14__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_14__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_15__CF_Inst_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_16__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_16__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_17__CF_Inst_n6,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_17__CF_Inst_n5,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_0__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_0__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_0__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_1__Compression1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_1__Compression2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_1__Compression3_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s1_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s2_n3,
         prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s3_n5,
         prince_rounds_AddKey1_forInv_XORInst_0_0_n3,
         prince_rounds_AddKey1_forInv_XORInst_0_1_n3,
         prince_rounds_AddKey1_forInv_XORInst_0_2_n3,
         prince_rounds_AddKey1_forInv_XORInst_0_3_n3,
         prince_rounds_AddKey1_forInv_XORInst_1_0_n3,
         prince_rounds_AddKey1_forInv_XORInst_1_1_n3,
         prince_rounds_AddKey1_forInv_XORInst_1_2_n3,
         prince_rounds_AddKey1_forInv_XORInst_1_3_n3,
         prince_rounds_AddKey1_forInv_XORInst_2_0_n3,
         prince_rounds_AddKey1_forInv_XORInst_2_1_n3,
         prince_rounds_AddKey1_forInv_XORInst_2_2_n3,
         prince_rounds_AddKey1_forInv_XORInst_2_3_n3,
         prince_rounds_AddKey1_forInv_XORInst_3_0_n3,
         prince_rounds_AddKey1_forInv_XORInst_3_1_n3,
         prince_rounds_AddKey1_forInv_XORInst_3_2_n3,
         prince_rounds_AddKey1_forInv_XORInst_3_3_n3,
         prince_rounds_AddKey1_forInv_XORInst_4_0_n3,
         prince_rounds_AddKey1_forInv_XORInst_4_1_n3,
         prince_rounds_AddKey1_forInv_XORInst_4_2_n3,
         prince_rounds_AddKey1_forInv_XORInst_4_3_n3,
         prince_rounds_AddKey1_forInv_XORInst_5_0_n3,
         prince_rounds_AddKey1_forInv_XORInst_5_1_n3,
         prince_rounds_AddKey1_forInv_XORInst_5_2_n3,
         prince_rounds_AddKey1_forInv_XORInst_5_3_n3,
         prince_rounds_AddKey1_forInv_XORInst_6_0_n3,
         prince_rounds_AddKey1_forInv_XORInst_6_1_n3,
         prince_rounds_AddKey1_forInv_XORInst_6_2_n3,
         prince_rounds_AddKey1_forInv_XORInst_6_3_n3,
         prince_rounds_AddKey1_forInv_XORInst_7_0_n3,
         prince_rounds_AddKey1_forInv_XORInst_7_1_n3,
         prince_rounds_AddKey1_forInv_XORInst_7_2_n3,
         prince_rounds_AddKey1_forInv_XORInst_7_3_n3,
         prince_rounds_AddKey1_forInv_XORInst_8_0_n3,
         prince_rounds_AddKey1_forInv_XORInst_8_1_n3,
         prince_rounds_AddKey1_forInv_XORInst_8_2_n3,
         prince_rounds_AddKey1_forInv_XORInst_8_3_n3,
         prince_rounds_AddKey1_forInv_XORInst_9_0_n3,
         prince_rounds_AddKey1_forInv_XORInst_9_1_n3,
         prince_rounds_AddKey1_forInv_XORInst_9_2_n3,
         prince_rounds_AddKey1_forInv_XORInst_9_3_n3,
         prince_rounds_AddKey1_forInv_XORInst_10_0_n3,
         prince_rounds_AddKey1_forInv_XORInst_10_1_n3,
         prince_rounds_AddKey1_forInv_XORInst_10_2_n3,
         prince_rounds_AddKey1_forInv_XORInst_10_3_n3,
         prince_rounds_AddKey1_forInv_XORInst_11_0_n3,
         prince_rounds_AddKey1_forInv_XORInst_11_1_n3,
         prince_rounds_AddKey1_forInv_XORInst_11_2_n3,
         prince_rounds_AddKey1_forInv_XORInst_11_3_n3,
         prince_rounds_AddKey1_forInv_XORInst_12_0_n3,
         prince_rounds_AddKey1_forInv_XORInst_12_1_n3,
         prince_rounds_AddKey1_forInv_XORInst_12_2_n3,
         prince_rounds_AddKey1_forInv_XORInst_12_3_n3,
         prince_rounds_AddKey1_forInv_XORInst_13_0_n3,
         prince_rounds_AddKey1_forInv_XORInst_13_1_n3,
         prince_rounds_AddKey1_forInv_XORInst_13_2_n3,
         prince_rounds_AddKey1_forInv_XORInst_13_3_n3,
         prince_rounds_AddKey1_forInv_XORInst_14_0_n3,
         prince_rounds_AddKey1_forInv_XORInst_14_1_n3,
         prince_rounds_AddKey1_forInv_XORInst_14_2_n3,
         prince_rounds_AddKey1_forInv_XORInst_14_3_n3,
         prince_rounds_AddKey1_forInv_XORInst_15_0_n3,
         prince_rounds_AddKey1_forInv_XORInst_15_1_n3,
         prince_rounds_AddKey1_forInv_XORInst_15_2_n3,
         prince_rounds_AddKey1_forInv_XORInst_15_3_n3,
         prince_rounds_AddKey2_forInv_XORInst_0_0_n3,
         prince_rounds_AddKey2_forInv_XORInst_0_1_n3,
         prince_rounds_AddKey2_forInv_XORInst_0_2_n3,
         prince_rounds_AddKey2_forInv_XORInst_0_3_n3,
         prince_rounds_AddKey2_forInv_XORInst_1_0_n3,
         prince_rounds_AddKey2_forInv_XORInst_1_1_n3,
         prince_rounds_AddKey2_forInv_XORInst_1_2_n3,
         prince_rounds_AddKey2_forInv_XORInst_1_3_n3,
         prince_rounds_AddKey2_forInv_XORInst_2_0_n3,
         prince_rounds_AddKey2_forInv_XORInst_2_1_n3,
         prince_rounds_AddKey2_forInv_XORInst_2_2_n3,
         prince_rounds_AddKey2_forInv_XORInst_2_3_n3,
         prince_rounds_AddKey2_forInv_XORInst_3_0_n3,
         prince_rounds_AddKey2_forInv_XORInst_3_1_n3,
         prince_rounds_AddKey2_forInv_XORInst_3_2_n3,
         prince_rounds_AddKey2_forInv_XORInst_3_3_n3,
         prince_rounds_AddKey2_forInv_XORInst_4_0_n3,
         prince_rounds_AddKey2_forInv_XORInst_4_1_n3,
         prince_rounds_AddKey2_forInv_XORInst_4_2_n3,
         prince_rounds_AddKey2_forInv_XORInst_4_3_n3,
         prince_rounds_AddKey2_forInv_XORInst_5_0_n3,
         prince_rounds_AddKey2_forInv_XORInst_5_1_n3,
         prince_rounds_AddKey2_forInv_XORInst_5_2_n3,
         prince_rounds_AddKey2_forInv_XORInst_5_3_n3,
         prince_rounds_AddKey2_forInv_XORInst_6_0_n3,
         prince_rounds_AddKey2_forInv_XORInst_6_1_n3,
         prince_rounds_AddKey2_forInv_XORInst_6_2_n3,
         prince_rounds_AddKey2_forInv_XORInst_6_3_n3,
         prince_rounds_AddKey2_forInv_XORInst_7_0_n3,
         prince_rounds_AddKey2_forInv_XORInst_7_1_n3,
         prince_rounds_AddKey2_forInv_XORInst_7_2_n3,
         prince_rounds_AddKey2_forInv_XORInst_7_3_n3,
         prince_rounds_AddKey2_forInv_XORInst_8_0_n3,
         prince_rounds_AddKey2_forInv_XORInst_8_1_n3,
         prince_rounds_AddKey2_forInv_XORInst_8_2_n3,
         prince_rounds_AddKey2_forInv_XORInst_8_3_n3,
         prince_rounds_AddKey2_forInv_XORInst_9_0_n3,
         prince_rounds_AddKey2_forInv_XORInst_9_1_n3,
         prince_rounds_AddKey2_forInv_XORInst_9_2_n3,
         prince_rounds_AddKey2_forInv_XORInst_9_3_n3,
         prince_rounds_AddKey2_forInv_XORInst_10_0_n3,
         prince_rounds_AddKey2_forInv_XORInst_10_1_n3,
         prince_rounds_AddKey2_forInv_XORInst_10_2_n3,
         prince_rounds_AddKey2_forInv_XORInst_10_3_n3,
         prince_rounds_AddKey2_forInv_XORInst_11_0_n3,
         prince_rounds_AddKey2_forInv_XORInst_11_1_n3,
         prince_rounds_AddKey2_forInv_XORInst_11_2_n3,
         prince_rounds_AddKey2_forInv_XORInst_11_3_n3,
         prince_rounds_AddKey2_forInv_XORInst_12_0_n3,
         prince_rounds_AddKey2_forInv_XORInst_12_1_n3,
         prince_rounds_AddKey2_forInv_XORInst_12_2_n3,
         prince_rounds_AddKey2_forInv_XORInst_12_3_n3,
         prince_rounds_AddKey2_forInv_XORInst_13_0_n3,
         prince_rounds_AddKey2_forInv_XORInst_13_1_n3,
         prince_rounds_AddKey2_forInv_XORInst_13_2_n3,
         prince_rounds_AddKey2_forInv_XORInst_13_3_n3,
         prince_rounds_AddKey2_forInv_XORInst_14_0_n3,
         prince_rounds_AddKey2_forInv_XORInst_14_1_n3,
         prince_rounds_AddKey2_forInv_XORInst_14_2_n3,
         prince_rounds_AddKey2_forInv_XORInst_14_3_n3,
         prince_rounds_AddKey2_forInv_XORInst_15_0_n3,
         prince_rounds_AddKey2_forInv_XORInst_15_1_n3,
         prince_rounds_AddKey2_forInv_XORInst_15_2_n3,
         prince_rounds_AddKey2_forInv_XORInst_15_3_n3,
         prince_rounds_AddKey3_forInv_XORInst_0_0_n3,
         prince_rounds_AddKey3_forInv_XORInst_0_1_n3,
         prince_rounds_AddKey3_forInv_XORInst_0_2_n3,
         prince_rounds_AddKey3_forInv_XORInst_0_3_n3,
         prince_rounds_AddKey3_forInv_XORInst_1_0_n3,
         prince_rounds_AddKey3_forInv_XORInst_1_1_n3,
         prince_rounds_AddKey3_forInv_XORInst_1_2_n3,
         prince_rounds_AddKey3_forInv_XORInst_1_3_n3,
         prince_rounds_AddKey3_forInv_XORInst_2_0_n3,
         prince_rounds_AddKey3_forInv_XORInst_2_1_n3,
         prince_rounds_AddKey3_forInv_XORInst_2_2_n3,
         prince_rounds_AddKey3_forInv_XORInst_2_3_n3,
         prince_rounds_AddKey3_forInv_XORInst_3_0_n3,
         prince_rounds_AddKey3_forInv_XORInst_3_1_n3,
         prince_rounds_AddKey3_forInv_XORInst_3_2_n3,
         prince_rounds_AddKey3_forInv_XORInst_3_3_n3,
         prince_rounds_AddKey3_forInv_XORInst_4_0_n3,
         prince_rounds_AddKey3_forInv_XORInst_4_1_n3,
         prince_rounds_AddKey3_forInv_XORInst_4_2_n3,
         prince_rounds_AddKey3_forInv_XORInst_4_3_n3,
         prince_rounds_AddKey3_forInv_XORInst_5_0_n3,
         prince_rounds_AddKey3_forInv_XORInst_5_1_n3,
         prince_rounds_AddKey3_forInv_XORInst_5_2_n3,
         prince_rounds_AddKey3_forInv_XORInst_5_3_n3,
         prince_rounds_AddKey3_forInv_XORInst_6_0_n3,
         prince_rounds_AddKey3_forInv_XORInst_6_1_n3,
         prince_rounds_AddKey3_forInv_XORInst_6_2_n3,
         prince_rounds_AddKey3_forInv_XORInst_6_3_n3,
         prince_rounds_AddKey3_forInv_XORInst_7_0_n3,
         prince_rounds_AddKey3_forInv_XORInst_7_1_n3,
         prince_rounds_AddKey3_forInv_XORInst_7_2_n3,
         prince_rounds_AddKey3_forInv_XORInst_7_3_n3,
         prince_rounds_AddKey3_forInv_XORInst_8_0_n3,
         prince_rounds_AddKey3_forInv_XORInst_8_1_n3,
         prince_rounds_AddKey3_forInv_XORInst_8_2_n3,
         prince_rounds_AddKey3_forInv_XORInst_8_3_n3,
         prince_rounds_AddKey3_forInv_XORInst_9_0_n3,
         prince_rounds_AddKey3_forInv_XORInst_9_1_n3,
         prince_rounds_AddKey3_forInv_XORInst_9_2_n3,
         prince_rounds_AddKey3_forInv_XORInst_9_3_n3,
         prince_rounds_AddKey3_forInv_XORInst_10_0_n3,
         prince_rounds_AddKey3_forInv_XORInst_10_1_n3,
         prince_rounds_AddKey3_forInv_XORInst_10_2_n3,
         prince_rounds_AddKey3_forInv_XORInst_10_3_n3,
         prince_rounds_AddKey3_forInv_XORInst_11_0_n3,
         prince_rounds_AddKey3_forInv_XORInst_11_1_n3,
         prince_rounds_AddKey3_forInv_XORInst_11_2_n3,
         prince_rounds_AddKey3_forInv_XORInst_11_3_n3,
         prince_rounds_AddKey3_forInv_XORInst_12_0_n3,
         prince_rounds_AddKey3_forInv_XORInst_12_1_n3,
         prince_rounds_AddKey3_forInv_XORInst_12_2_n3,
         prince_rounds_AddKey3_forInv_XORInst_12_3_n3,
         prince_rounds_AddKey3_forInv_XORInst_13_0_n3,
         prince_rounds_AddKey3_forInv_XORInst_13_1_n3,
         prince_rounds_AddKey3_forInv_XORInst_13_2_n3,
         prince_rounds_AddKey3_forInv_XORInst_13_3_n3,
         prince_rounds_AddKey3_forInv_XORInst_14_0_n3,
         prince_rounds_AddKey3_forInv_XORInst_14_1_n3,
         prince_rounds_AddKey3_forInv_XORInst_14_2_n3,
         prince_rounds_AddKey3_forInv_XORInst_14_3_n3,
         prince_rounds_AddKey3_forInv_XORInst_15_0_n3,
         prince_rounds_AddKey3_forInv_XORInst_15_1_n3,
         prince_rounds_AddKey3_forInv_XORInst_15_2_n3,
         prince_rounds_AddKey3_forInv_XORInst_15_3_n3,
         prince_rounds_S_Sinv_mul1_n10, prince_rounds_S_Sinv_mul1_n9,
         prince_rounds_S_Sinv_mul1_n8, prince_rounds_S_Sinv_mul1_n7,
         prince_rounds_S_Sinv_mul2_n10, prince_rounds_S_Sinv_mul2_n9,
         prince_rounds_S_Sinv_mul2_n8, prince_rounds_S_Sinv_mul2_n7,
         prince_rounds_S_Sinv_mul3_n8, prince_rounds_S_Sinv_mul3_n7,
         prince_rounds_S_Sinv_mul3_n6, prince_rounds_mul_s1_n96,
         prince_rounds_mul_s1_n95, prince_rounds_mul_s1_n94,
         prince_rounds_mul_s1_n93, prince_rounds_mul_s1_n92,
         prince_rounds_mul_s1_n91, prince_rounds_mul_s1_n90,
         prince_rounds_mul_s1_n89, prince_rounds_mul_s1_n88,
         prince_rounds_mul_s1_n87, prince_rounds_mul_s1_n86,
         prince_rounds_mul_s1_n85, prince_rounds_mul_s1_n84,
         prince_rounds_mul_s1_n83, prince_rounds_mul_s1_n82,
         prince_rounds_mul_s1_n81, prince_rounds_mul_s1_n80,
         prince_rounds_mul_s1_n79, prince_rounds_mul_s1_n78,
         prince_rounds_mul_s1_n77, prince_rounds_mul_s1_n76,
         prince_rounds_mul_s1_n75, prince_rounds_mul_s1_n74,
         prince_rounds_mul_s1_n73, prince_rounds_mul_s1_n72,
         prince_rounds_mul_s1_n71, prince_rounds_mul_s1_n70,
         prince_rounds_mul_s1_n69, prince_rounds_mul_s1_n68,
         prince_rounds_mul_s1_n67, prince_rounds_mul_s1_n66,
         prince_rounds_mul_s1_n65, prince_rounds_mul_s2_n96,
         prince_rounds_mul_s2_n95, prince_rounds_mul_s2_n94,
         prince_rounds_mul_s2_n93, prince_rounds_mul_s2_n92,
         prince_rounds_mul_s2_n91, prince_rounds_mul_s2_n90,
         prince_rounds_mul_s2_n89, prince_rounds_mul_s2_n88,
         prince_rounds_mul_s2_n87, prince_rounds_mul_s2_n86,
         prince_rounds_mul_s2_n85, prince_rounds_mul_s2_n84,
         prince_rounds_mul_s2_n83, prince_rounds_mul_s2_n82,
         prince_rounds_mul_s2_n81, prince_rounds_mul_s2_n80,
         prince_rounds_mul_s2_n79, prince_rounds_mul_s2_n78,
         prince_rounds_mul_s2_n77, prince_rounds_mul_s2_n76,
         prince_rounds_mul_s2_n75, prince_rounds_mul_s2_n74,
         prince_rounds_mul_s2_n73, prince_rounds_mul_s2_n72,
         prince_rounds_mul_s2_n71, prince_rounds_mul_s2_n70,
         prince_rounds_mul_s2_n69, prince_rounds_mul_s2_n68,
         prince_rounds_mul_s2_n67, prince_rounds_mul_s2_n66,
         prince_rounds_mul_s2_n65, prince_rounds_mul_s3_n96,
         prince_rounds_mul_s3_n95, prince_rounds_mul_s3_n94,
         prince_rounds_mul_s3_n93, prince_rounds_mul_s3_n92,
         prince_rounds_mul_s3_n91, prince_rounds_mul_s3_n90,
         prince_rounds_mul_s3_n89, prince_rounds_mul_s3_n88,
         prince_rounds_mul_s3_n87, prince_rounds_mul_s3_n86,
         prince_rounds_mul_s3_n85, prince_rounds_mul_s3_n84,
         prince_rounds_mul_s3_n83, prince_rounds_mul_s3_n82,
         prince_rounds_mul_s3_n81, prince_rounds_mul_s3_n80,
         prince_rounds_mul_s3_n79, prince_rounds_mul_s3_n78,
         prince_rounds_mul_s3_n77, prince_rounds_mul_s3_n76,
         prince_rounds_mul_s3_n75, prince_rounds_mul_s3_n74,
         prince_rounds_mul_s3_n73, prince_rounds_mul_s3_n72,
         prince_rounds_mul_s3_n71, prince_rounds_mul_s3_n70,
         prince_rounds_mul_s3_n69, prince_rounds_mul_s3_n68,
         prince_rounds_mul_s3_n67, prince_rounds_mul_s3_n66,
         prince_rounds_mul_s3_n65, prince_AddKeyOut1_XORInst_0_0_n3,
         prince_AddKeyOut1_XORInst_0_1_n3, prince_AddKeyOut1_XORInst_0_2_n3,
         prince_AddKeyOut1_XORInst_0_3_n3, prince_AddKeyOut1_XORInst_1_0_n3,
         prince_AddKeyOut1_XORInst_1_1_n3, prince_AddKeyOut1_XORInst_1_2_n3,
         prince_AddKeyOut1_XORInst_1_3_n3, prince_AddKeyOut1_XORInst_2_0_n3,
         prince_AddKeyOut1_XORInst_2_1_n3, prince_AddKeyOut1_XORInst_2_2_n3,
         prince_AddKeyOut1_XORInst_2_3_n3, prince_AddKeyOut1_XORInst_3_0_n3,
         prince_AddKeyOut1_XORInst_3_1_n3, prince_AddKeyOut1_XORInst_3_2_n3,
         prince_AddKeyOut1_XORInst_3_3_n3, prince_AddKeyOut1_XORInst_4_0_n3,
         prince_AddKeyOut1_XORInst_4_1_n3, prince_AddKeyOut1_XORInst_4_2_n3,
         prince_AddKeyOut1_XORInst_4_3_n3, prince_AddKeyOut1_XORInst_5_0_n3,
         prince_AddKeyOut1_XORInst_5_1_n3, prince_AddKeyOut1_XORInst_5_2_n3,
         prince_AddKeyOut1_XORInst_5_3_n3, prince_AddKeyOut1_XORInst_6_0_n3,
         prince_AddKeyOut1_XORInst_6_1_n3, prince_AddKeyOut1_XORInst_6_2_n3,
         prince_AddKeyOut1_XORInst_6_3_n3, prince_AddKeyOut1_XORInst_7_0_n3,
         prince_AddKeyOut1_XORInst_7_1_n3, prince_AddKeyOut1_XORInst_7_2_n3,
         prince_AddKeyOut1_XORInst_7_3_n3, prince_AddKeyOut1_XORInst_8_0_n3,
         prince_AddKeyOut1_XORInst_8_1_n3, prince_AddKeyOut1_XORInst_8_2_n3,
         prince_AddKeyOut1_XORInst_8_3_n3, prince_AddKeyOut1_XORInst_9_0_n3,
         prince_AddKeyOut1_XORInst_9_1_n3, prince_AddKeyOut1_XORInst_9_2_n3,
         prince_AddKeyOut1_XORInst_9_3_n3, prince_AddKeyOut1_XORInst_10_0_n3,
         prince_AddKeyOut1_XORInst_10_1_n3, prince_AddKeyOut1_XORInst_10_2_n3,
         prince_AddKeyOut1_XORInst_10_3_n3, prince_AddKeyOut1_XORInst_11_0_n3,
         prince_AddKeyOut1_XORInst_11_1_n3, prince_AddKeyOut1_XORInst_11_2_n3,
         prince_AddKeyOut1_XORInst_11_3_n3, prince_AddKeyOut1_XORInst_12_0_n3,
         prince_AddKeyOut1_XORInst_12_1_n3, prince_AddKeyOut1_XORInst_12_2_n3,
         prince_AddKeyOut1_XORInst_12_3_n3, prince_AddKeyOut1_XORInst_13_0_n3,
         prince_AddKeyOut1_XORInst_13_1_n3, prince_AddKeyOut1_XORInst_13_2_n3,
         prince_AddKeyOut1_XORInst_13_3_n3, prince_AddKeyOut1_XORInst_14_0_n3,
         prince_AddKeyOut1_XORInst_14_1_n3, prince_AddKeyOut1_XORInst_14_2_n3,
         prince_AddKeyOut1_XORInst_14_3_n3, prince_AddKeyOut1_XORInst_15_0_n3,
         prince_AddKeyOut1_XORInst_15_1_n3, prince_AddKeyOut1_XORInst_15_2_n3,
         prince_AddKeyOut1_XORInst_15_3_n3, prince_AddKeyOut2_XORInst_0_0_n3,
         prince_AddKeyOut2_XORInst_0_1_n3, prince_AddKeyOut2_XORInst_0_2_n3,
         prince_AddKeyOut2_XORInst_0_3_n3, prince_AddKeyOut2_XORInst_1_0_n3,
         prince_AddKeyOut2_XORInst_1_1_n3, prince_AddKeyOut2_XORInst_1_2_n3,
         prince_AddKeyOut2_XORInst_1_3_n3, prince_AddKeyOut2_XORInst_2_0_n3,
         prince_AddKeyOut2_XORInst_2_1_n3, prince_AddKeyOut2_XORInst_2_2_n3,
         prince_AddKeyOut2_XORInst_2_3_n3, prince_AddKeyOut2_XORInst_3_0_n3,
         prince_AddKeyOut2_XORInst_3_1_n3, prince_AddKeyOut2_XORInst_3_2_n3,
         prince_AddKeyOut2_XORInst_3_3_n3, prince_AddKeyOut2_XORInst_4_0_n3,
         prince_AddKeyOut2_XORInst_4_1_n3, prince_AddKeyOut2_XORInst_4_2_n3,
         prince_AddKeyOut2_XORInst_4_3_n3, prince_AddKeyOut2_XORInst_5_0_n3,
         prince_AddKeyOut2_XORInst_5_1_n3, prince_AddKeyOut2_XORInst_5_2_n3,
         prince_AddKeyOut2_XORInst_5_3_n3, prince_AddKeyOut2_XORInst_6_0_n3,
         prince_AddKeyOut2_XORInst_6_1_n3, prince_AddKeyOut2_XORInst_6_2_n3,
         prince_AddKeyOut2_XORInst_6_3_n3, prince_AddKeyOut2_XORInst_7_0_n3,
         prince_AddKeyOut2_XORInst_7_1_n3, prince_AddKeyOut2_XORInst_7_2_n3,
         prince_AddKeyOut2_XORInst_7_3_n3, prince_AddKeyOut2_XORInst_8_0_n3,
         prince_AddKeyOut2_XORInst_8_1_n3, prince_AddKeyOut2_XORInst_8_2_n3,
         prince_AddKeyOut2_XORInst_8_3_n3, prince_AddKeyOut2_XORInst_9_0_n3,
         prince_AddKeyOut2_XORInst_9_1_n3, prince_AddKeyOut2_XORInst_9_2_n3,
         prince_AddKeyOut2_XORInst_9_3_n3, prince_AddKeyOut2_XORInst_10_0_n3,
         prince_AddKeyOut2_XORInst_10_1_n3, prince_AddKeyOut2_XORInst_10_2_n3,
         prince_AddKeyOut2_XORInst_10_3_n3, prince_AddKeyOut2_XORInst_11_0_n3,
         prince_AddKeyOut2_XORInst_11_1_n3, prince_AddKeyOut2_XORInst_11_2_n3,
         prince_AddKeyOut2_XORInst_11_3_n3, prince_AddKeyOut2_XORInst_12_0_n3,
         prince_AddKeyOut2_XORInst_12_1_n3, prince_AddKeyOut2_XORInst_12_2_n3,
         prince_AddKeyOut2_XORInst_12_3_n3, prince_AddKeyOut2_XORInst_13_0_n3,
         prince_AddKeyOut2_XORInst_13_1_n3, prince_AddKeyOut2_XORInst_13_2_n3,
         prince_AddKeyOut2_XORInst_13_3_n3, prince_AddKeyOut2_XORInst_14_0_n3,
         prince_AddKeyOut2_XORInst_14_1_n3, prince_AddKeyOut2_XORInst_14_2_n3,
         prince_AddKeyOut2_XORInst_14_3_n3, prince_AddKeyOut2_XORInst_15_0_n3,
         prince_AddKeyOut2_XORInst_15_1_n3, prince_AddKeyOut2_XORInst_15_2_n3,
         prince_AddKeyOut2_XORInst_15_3_n3, prince_AddKeyOut3_XORInst_0_0_n3,
         prince_AddKeyOut3_XORInst_0_1_n3, prince_AddKeyOut3_XORInst_0_2_n3,
         prince_AddKeyOut3_XORInst_0_3_n3, prince_AddKeyOut3_XORInst_1_0_n3,
         prince_AddKeyOut3_XORInst_1_1_n3, prince_AddKeyOut3_XORInst_1_2_n3,
         prince_AddKeyOut3_XORInst_1_3_n3, prince_AddKeyOut3_XORInst_2_0_n3,
         prince_AddKeyOut3_XORInst_2_1_n3, prince_AddKeyOut3_XORInst_2_2_n3,
         prince_AddKeyOut3_XORInst_2_3_n3, prince_AddKeyOut3_XORInst_3_0_n3,
         prince_AddKeyOut3_XORInst_3_1_n3, prince_AddKeyOut3_XORInst_3_2_n3,
         prince_AddKeyOut3_XORInst_3_3_n3, prince_AddKeyOut3_XORInst_4_0_n3,
         prince_AddKeyOut3_XORInst_4_1_n3, prince_AddKeyOut3_XORInst_4_2_n3,
         prince_AddKeyOut3_XORInst_4_3_n3, prince_AddKeyOut3_XORInst_5_0_n3,
         prince_AddKeyOut3_XORInst_5_1_n3, prince_AddKeyOut3_XORInst_5_2_n3,
         prince_AddKeyOut3_XORInst_5_3_n3, prince_AddKeyOut3_XORInst_6_0_n3,
         prince_AddKeyOut3_XORInst_6_1_n3, prince_AddKeyOut3_XORInst_6_2_n3,
         prince_AddKeyOut3_XORInst_6_3_n3, prince_AddKeyOut3_XORInst_7_0_n3,
         prince_AddKeyOut3_XORInst_7_1_n3, prince_AddKeyOut3_XORInst_7_2_n3,
         prince_AddKeyOut3_XORInst_7_3_n3, prince_AddKeyOut3_XORInst_8_0_n3,
         prince_AddKeyOut3_XORInst_8_1_n3, prince_AddKeyOut3_XORInst_8_2_n3,
         prince_AddKeyOut3_XORInst_8_3_n3, prince_AddKeyOut3_XORInst_9_0_n3,
         prince_AddKeyOut3_XORInst_9_1_n3, prince_AddKeyOut3_XORInst_9_2_n3,
         prince_AddKeyOut3_XORInst_9_3_n3, prince_AddKeyOut3_XORInst_10_0_n3,
         prince_AddKeyOut3_XORInst_10_1_n3, prince_AddKeyOut3_XORInst_10_2_n3,
         prince_AddKeyOut3_XORInst_10_3_n3, prince_AddKeyOut3_XORInst_11_0_n3,
         prince_AddKeyOut3_XORInst_11_1_n3, prince_AddKeyOut3_XORInst_11_2_n3,
         prince_AddKeyOut3_XORInst_11_3_n3, prince_AddKeyOut3_XORInst_12_0_n3,
         prince_AddKeyOut3_XORInst_12_1_n3, prince_AddKeyOut3_XORInst_12_2_n3,
         prince_AddKeyOut3_XORInst_12_3_n3, prince_AddKeyOut3_XORInst_13_0_n3,
         prince_AddKeyOut3_XORInst_13_1_n3, prince_AddKeyOut3_XORInst_13_2_n3,
         prince_AddKeyOut3_XORInst_13_3_n3, prince_AddKeyOut3_XORInst_14_0_n3,
         prince_AddKeyOut3_XORInst_14_1_n3, prince_AddKeyOut3_XORInst_14_2_n3,
         prince_AddKeyOut3_XORInst_14_3_n3, prince_AddKeyOut3_XORInst_15_0_n3,
         prince_AddKeyOut3_XORInst_15_1_n3, prince_AddKeyOut3_XORInst_15_2_n3,
         prince_AddKeyOut3_XORInst_15_3_n3;
  wire   [3:0] round_Signal;
  wire   [63:0] prince_rounds_Output_s3;
  wire   [63:0] prince_rounds_Output_s2;
  wire   [63:0] prince_rounds_Output_s1;
  wire   [63:0] prince_SR_Inv_Result_s3;
  wire   [63:0] prince_SR_Inv_Result_s2;
  wire   [63:0] prince_SR_Inv_Result_s1;
  wire   [63:0] prince_rounds_mul_input_s3;
  wire   [63:0] prince_rounds_mul_input_s2;
  wire   [63:0] prince_rounds_mul_input_s1;
  wire   [63:0] prince_rounds_SR_Inv_Result_s3;
  wire   [63:0] prince_rounds_SR_Inv_Result_s2;
  wire   [63:0] prince_rounds_SR_Inv_Result_s1;
  wire   [62:0] prince_rounds_sub_Inv_Result_s3;
  wire   [61:1] prince_rounds_sub_Inv_Result_s2;
  wire   [61:1] prince_rounds_sub_Inv_Result_s1;
  wire   [63:0] prince_rounds_sub_Result_s3;
  wire   [63:0] prince_rounds_sub_Result_s2;
  wire   [63:0] prince_rounds_sub_Result_s1;
  wire   [63:0] prince_rounds_round_inputXORkeyRCON_s3;
  wire   [63:0] prince_rounds_round_inputXORkeyRCON_s2;
  wire   [63:0] prince_rounds_round_inputXORkeyRCON_s1;
  wire   [63:0] prince_rounds_SR_Result_s3;
  wire   [63:0] prince_rounds_SR_Result_s2;
  wire   [63:0] prince_rounds_SR_Result_s1;
  wire   [63:0] prince_rounds_mul_result_s3;
  wire   [63:0] prince_rounds_mul_result_s2;
  wire   [63:0] prince_rounds_mul_result_s1;
  wire   [63:1] prince_rounds_round_Constant;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_2_out1;
  wire   [1:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_2_out1;
  wire   [1:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_2_out1;
  wire   [1:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_2_out1;
  wire   [1:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_2_out1;
  wire   [1:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_2_out1;
  wire   [1:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_2_out1;
  wire   [1:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_2_out1;
  wire   [1:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_2_out1;
  wire   [1:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_2_out1;
  wire   [1:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_2_out1;
  wire   [1:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out
;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_2_out1;
  wire   [1:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out
;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_2_out1;
  wire   [1:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out
;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_2_out1;
  wire   [1:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out
;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_2_out1;
  wire   [1:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out
;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_2_out1;
  wire   [1:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2;
  wire   [3:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg
;
  wire   [17:0] prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out
;

  AOI22_X1 MyController_U45 ( .A1(MyController_n36), .A2(MyController_n38), 
        .B1(MyController_n35), .B2(MyController_n34), .ZN(MyController_n77) );
  AOI22_X1 MyController_U44 ( .A1(MyController_n36), .A2(MyController_n8), 
        .B1(MyController_n33), .B2(MyController_n34), .ZN(MyController_n76) );
  INV_X1 MyController_U43 ( .A(MyController_n36), .ZN(MyController_n34) );
  MUX2_X1 MyController_U42 ( .A(round_Signal[2]), .B(MyController_n43), .S(
        MyController_n36), .Z(MyController_n75) );
  NOR2_X1 MyController_U41 ( .A1(reset), .A2(MyController_n32), .ZN(
        MyController_n36) );
  AOI211_X1 MyController_U40 ( .C1(MyController_n31), .C2(MyController_n6), 
        .A(reset), .B(MyController_n29), .ZN(round_Signal[2]) );
  AOI21_X1 MyController_U39 ( .B1(MyController_n30), .B2(MyController_n28), 
        .A(MyController_n27), .ZN(MyController_n74) );
  OAI21_X1 MyController_U38 ( .B1(MyController_n30), .B2(MyController_n28), 
        .A(MyController_n10), .ZN(MyController_n27) );
  NAND4_X1 MyController_U37 ( .A1(MyController_n40), .A2(MyController_n26), 
        .A3(MyController_n29), .A4(MyController_n9), .ZN(MyController_n28) );
  NOR4_X1 MyController_U36 ( .A1(MyController_n6), .A2(MyController_n25), .A3(
        round_Signal[1]), .A4(MyController_n35), .ZN(done) );
  INV_X1 MyController_U35 ( .A(round_Signal[0]), .ZN(MyController_n35) );
  OR2_X1 MyController_U34 ( .A1(round_Signal[3]), .A2(MyController_n19), .ZN(
        MyController_N25) );
  AND2_X1 MyController_U33 ( .A1(MyController_n23), .A2(MyController_n18), 
        .ZN(MyController_N19) );
  NOR3_X1 MyController_U32 ( .A1(MyController_n17), .A2(MyController_n22), 
        .A3(MyController_n32), .ZN(MyController_N18) );
  NOR2_X1 MyController_U31 ( .A1(MyController_n20), .A2(MyController_n16), 
        .ZN(MyController_n22) );
  AOI211_X1 MyController_U30 ( .C1(MyController_n4), .C2(MyController_n21), 
        .A(MyController_n20), .B(MyController_n32), .ZN(MyController_N17) );
  OAI21_X1 MyController_U29 ( .B1(MyController_n15), .B2(MyController_n23), 
        .A(MyController_n18), .ZN(MyController_n32) );
  NAND2_X1 MyController_U28 ( .A1(MyController_n19), .A2(MyController_n25), 
        .ZN(MyController_n18) );
  INV_X1 MyController_U27 ( .A(round_Signal[3]), .ZN(MyController_n25) );
  NOR4_X1 MyController_U26 ( .A1(MyController_n14), .A2(MyController_n13), 
        .A3(MyController_n16), .A4(MyController_n24), .ZN(MyController_n19) );
  INV_X1 MyController_U25 ( .A(MyController_n20), .ZN(MyController_n13) );
  INV_X1 MyController_U24 ( .A(MyController_n14), .ZN(MyController_n23) );
  XNOR2_X1 MyController_U23 ( .A(MyController_n12), .B(MyController_n17), .ZN(
        MyController_n14) );
  AND2_X1 MyController_U22 ( .A1(MyController_n20), .A2(MyController_n16), 
        .ZN(MyController_n17) );
  NAND2_X1 MyController_U21 ( .A1(MyController_n47), .A2(MyController_n10), 
        .ZN(MyController_n16) );
  NAND2_X1 MyController_U20 ( .A1(MyController_n40), .A2(MyController_n10), 
        .ZN(MyController_n12) );
  OAI211_X1 MyController_U19 ( .C1(round_Signal[3]), .C2(MyController_n24), 
        .A(MyController_n26), .B(MyController_n21), .ZN(MyController_n15) );
  NOR2_X1 MyController_U18 ( .A1(MyController_n47), .A2(MyController_n44), 
        .ZN(MyController_n26) );
  NAND3_X1 MyController_U17 ( .A1(MyController_n43), .A2(round_Signal[0]), 
        .A3(round_Signal[1]), .ZN(MyController_n24) );
  AOI221_X1 MyController_U16 ( .B1(MyController_n30), .B2(MyController_n11), 
        .C1(MyController_n7), .C2(MyController_n29), .A(reset), .ZN(
        round_Signal[3]) );
  INV_X1 MyController_U15 ( .A(MyController_n29), .ZN(MyController_n11) );
  NOR2_X1 MyController_U14 ( .A1(MyController_n31), .A2(MyController_n6), .ZN(
        MyController_n29) );
  NOR2_X1 MyController_U13 ( .A1(MyController_n21), .A2(MyController_n4), .ZN(
        MyController_n20) );
  NOR2_X1 MyController_U12 ( .A1(reset), .A2(MyController_n46), .ZN(
        MyController_n21) );
  NOR2_X1 MyController_U11 ( .A1(reset), .A2(MyController_n5), .ZN(
        round_Signal[0]) );
  INV_X1 MyController_U10 ( .A(MyController_n33), .ZN(round_Signal[1]) );
  AOI221_X1 MyController_U9 ( .B1(MyController_n31), .B2(MyController_n5), 
        .C1(MyController_n31), .C2(MyController_n45), .A(reset), .ZN(
        MyController_n33) );
  NAND2_X1 MyController_U8 ( .A1(MyController_n5), .A2(MyController_n45), .ZN(
        MyController_n31) );
  INV_X1 MyController_U7 ( .A(reset), .ZN(MyController_n10) );
  AND2_X1 MyController_U6 ( .A1(MyController_n10), .A2(MyController_n44), .ZN(
        MyController_n4) );
  OAI21_X1 MyController_U5 ( .B1(MyController_n24), .B2(MyController_n3), .A(
        MyController_n25), .ZN(MyController_N27) );
  NOR2_X1 MyController_U4 ( .A1(MyController_n23), .A2(MyController_n2), .ZN(
        MyController_n3) );
  AOI211_X1 MyController_U3 ( .C1(MyController_n21), .C2(MyController_n4), .A(
        MyController_n20), .B(MyController_n22), .ZN(MyController_n2) );
  DFF_X1 MyController_roundEnd_Select_reg ( .D(MyController_N25), .CK(clk), 
        .Q(roundEnd_Select_Signal), .QN() );
  DFF_X1 MyController_roundHalf_Select_reg ( .D(MyController_N27), .CK(clk), 
        .Q(roundHalf_Select_Signal), .QN() );
  DFF_X1 MyController_RoundCounterReg_reg_3_ ( .D(MyController_n74), .CK(clk), 
        .Q(MyController_n7), .QN(MyController_n30) );
  DFF_X1 MyController_PerRoundCounterReg_reg_1_ ( .D(MyController_N17), .CK(
        clk), .Q(MyController_n46), .QN(MyController_n9) );
  DFF_X1 MyController_PerRoundCounterReg_reg_2_ ( .D(MyController_N18), .CK(
        clk), .Q(), .QN(MyController_n47) );
  DFF_X1 MyController_PerRoundCounterReg_reg_3_ ( .D(MyController_N19), .CK(
        clk), .Q(), .QN(MyController_n40) );
  DFF_X1 MyController_RoundCounterReg_reg_2_ ( .D(MyController_n75), .CK(clk), 
        .Q(MyController_n43), .QN(MyController_n6) );
  DFF_X1 MyController_RoundCounterReg_reg_1_ ( .D(MyController_n76), .CK(clk), 
        .Q(MyController_n45), .QN(MyController_n8) );
  DFF_X1 MyController_RoundCounterReg_reg_0_ ( .D(MyController_n77), .CK(clk), 
        .Q(MyController_n5), .QN(MyController_n38) );
  DFF_X1 MyController_PerRoundCounterReg_reg_0_ ( .D(MyController_n4), .CK(clk), .Q(), .QN(MyController_n44) );
  XOR2_X1 prince_U3 ( .A(enc_dec), .B(reset), .Z(prince_enc_dec_xor_reset) );
  BUF_X1 prince_U2 ( .A(prince_enc_dec_xor_reset), .Z(prince_n3) );
  XOR2_X1 prince_KeyDriv1_U1 ( .A(Key1[127]), .B(Key1[65]), .Z(
        prince_k_0_p_share1_0_) );
  XOR2_X1 prince_KeyDriv2_U1 ( .A(Key2[127]), .B(Key2[65]), .Z(
        prince_k_0_p_share2_0_) );
  XOR2_X1 prince_KeyDriv3_U1 ( .A(Key3[127]), .B(Key3[65]), .Z(
        prince_k_0_p_share3_0_) );
  BUF_X1 prince_KeyMUX1_U4 ( .A(prince_n3), .Z(prince_KeyMUX1_n7) );
  BUF_X1 prince_KeyMUX1_U3 ( .A(prince_KeyMUX1_n7), .Z(prince_KeyMUX1_n9) );
  BUF_X1 prince_KeyMUX1_U2 ( .A(prince_n3), .Z(prince_KeyMUX1_n8) );
  BUF_X1 prince_KeyMUX1_U1 ( .A(prince_KeyMUX1_n8), .Z(prince_KeyMUX1_n10) );
  MUX2_X1 prince_KeyMUX1_MUXInst_0_U1 ( .A(prince_k_0_p_share1_0_), .B(
        Key1[64]), .S(prince_KeyMUX1_n8), .Z(prince_selected_Key1_0_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_1_U1 ( .A(Key1[66]), .B(Key1[65]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_1_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_2_U1 ( .A(Key1[67]), .B(Key1[66]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_2_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_3_U1 ( .A(Key1[68]), .B(Key1[67]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_3_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_4_U1 ( .A(Key1[69]), .B(Key1[68]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_4_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_5_U1 ( .A(Key1[70]), .B(Key1[69]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_5_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_6_U1 ( .A(Key1[71]), .B(Key1[70]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_6_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_7_U1 ( .A(Key1[72]), .B(Key1[71]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_7_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_8_U1 ( .A(Key1[73]), .B(Key1[72]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_8_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_9_U1 ( .A(Key1[74]), .B(Key1[73]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_9_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_10_U1 ( .A(Key1[75]), .B(Key1[74]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_10_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_11_U1 ( .A(Key1[76]), .B(Key1[75]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_11_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_12_U1 ( .A(Key1[77]), .B(Key1[76]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_12_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_13_U1 ( .A(Key1[78]), .B(Key1[77]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_13_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_14_U1 ( .A(Key1[79]), .B(Key1[78]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_14_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_15_U1 ( .A(Key1[80]), .B(Key1[79]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_15_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_16_U1 ( .A(Key1[81]), .B(Key1[80]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_16_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_17_U1 ( .A(Key1[82]), .B(Key1[81]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_17_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_18_U1 ( .A(Key1[83]), .B(Key1[82]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_18_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_19_U1 ( .A(Key1[84]), .B(Key1[83]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_19_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_20_U1 ( .A(Key1[85]), .B(Key1[84]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_20_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_21_U1 ( .A(Key1[86]), .B(Key1[85]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_21_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_22_U1 ( .A(Key1[87]), .B(Key1[86]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_22_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_23_U1 ( .A(Key1[88]), .B(Key1[87]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_23_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_24_U1 ( .A(Key1[89]), .B(Key1[88]), .S(
        prince_KeyMUX1_n7), .Z(prince_selected_Key1_24_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_25_U1 ( .A(Key1[90]), .B(Key1[89]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_25_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_26_U1 ( .A(Key1[91]), .B(Key1[90]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_26_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_27_U1 ( .A(Key1[92]), .B(Key1[91]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_27_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_28_U1 ( .A(Key1[93]), .B(Key1[92]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_28_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_29_U1 ( .A(Key1[94]), .B(Key1[93]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_29_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_30_U1 ( .A(Key1[95]), .B(Key1[94]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_30_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_31_U1 ( .A(Key1[96]), .B(Key1[95]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_31_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_32_U1 ( .A(Key1[97]), .B(Key1[96]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_32_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_33_U1 ( .A(Key1[98]), .B(Key1[97]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_33_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_34_U1 ( .A(Key1[99]), .B(Key1[98]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_34_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_35_U1 ( .A(Key1[100]), .B(Key1[99]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_35_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_36_U1 ( .A(Key1[101]), .B(Key1[100]), .S(
        prince_KeyMUX1_n9), .Z(prince_selected_Key1_36_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_37_U1 ( .A(Key1[102]), .B(Key1[101]), .S(
        prince_KeyMUX1_n10), .Z(prince_selected_Key1_37_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_38_U1 ( .A(Key1[103]), .B(Key1[102]), .S(
        prince_KeyMUX1_n8), .Z(prince_selected_Key1_38_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_39_U1 ( .A(Key1[104]), .B(Key1[103]), .S(
        prince_KeyMUX1_n10), .Z(prince_selected_Key1_39_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_40_U1 ( .A(Key1[105]), .B(Key1[104]), .S(
        prince_KeyMUX1_n8), .Z(prince_selected_Key1_40_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_41_U1 ( .A(Key1[106]), .B(Key1[105]), .S(
        prince_KeyMUX1_n10), .Z(prince_selected_Key1_41_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_42_U1 ( .A(Key1[107]), .B(Key1[106]), .S(
        prince_KeyMUX1_n8), .Z(prince_selected_Key1_42_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_43_U1 ( .A(Key1[108]), .B(Key1[107]), .S(
        prince_KeyMUX1_n8), .Z(prince_selected_Key1_43_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_44_U1 ( .A(Key1[109]), .B(Key1[108]), .S(
        prince_KeyMUX1_n8), .Z(prince_selected_Key1_44_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_45_U1 ( .A(Key1[110]), .B(Key1[109]), .S(
        prince_KeyMUX1_n8), .Z(prince_selected_Key1_45_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_46_U1 ( .A(Key1[111]), .B(Key1[110]), .S(
        prince_KeyMUX1_n8), .Z(prince_selected_Key1_46_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_47_U1 ( .A(Key1[112]), .B(Key1[111]), .S(
        prince_KeyMUX1_n8), .Z(prince_selected_Key1_47_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_48_U1 ( .A(Key1[113]), .B(Key1[112]), .S(
        prince_KeyMUX1_n8), .Z(prince_selected_Key1_48_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_49_U1 ( .A(Key1[114]), .B(Key1[113]), .S(
        prince_KeyMUX1_n10), .Z(prince_selected_Key1_49_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_50_U1 ( .A(Key1[115]), .B(Key1[114]), .S(
        prince_KeyMUX1_n10), .Z(prince_selected_Key1_50_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_51_U1 ( .A(Key1[116]), .B(Key1[115]), .S(
        prince_KeyMUX1_n10), .Z(prince_selected_Key1_51_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_52_U1 ( .A(Key1[117]), .B(Key1[116]), .S(
        prince_KeyMUX1_n10), .Z(prince_selected_Key1_52_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_53_U1 ( .A(Key1[118]), .B(Key1[117]), .S(
        prince_KeyMUX1_n10), .Z(prince_selected_Key1_53_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_54_U1 ( .A(Key1[119]), .B(Key1[118]), .S(
        prince_KeyMUX1_n10), .Z(prince_selected_Key1_54_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_55_U1 ( .A(Key1[120]), .B(Key1[119]), .S(
        prince_KeyMUX1_n10), .Z(prince_selected_Key1_55_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_56_U1 ( .A(Key1[121]), .B(Key1[120]), .S(
        prince_KeyMUX1_n10), .Z(prince_selected_Key1_56_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_57_U1 ( .A(Key1[122]), .B(Key1[121]), .S(
        prince_KeyMUX1_n10), .Z(prince_selected_Key1_57_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_58_U1 ( .A(Key1[123]), .B(Key1[122]), .S(
        prince_KeyMUX1_n10), .Z(prince_selected_Key1_58_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_59_U1 ( .A(Key1[124]), .B(Key1[123]), .S(
        prince_KeyMUX1_n10), .Z(prince_selected_Key1_59_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_60_U1 ( .A(Key1[125]), .B(Key1[124]), .S(
        prince_KeyMUX1_n10), .Z(prince_selected_Key1_60_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_61_U1 ( .A(Key1[126]), .B(Key1[125]), .S(
        prince_KeyMUX1_n8), .Z(prince_selected_Key1_61_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_62_U1 ( .A(Key1[127]), .B(Key1[126]), .S(
        prince_KeyMUX1_n8), .Z(prince_selected_Key1_62_) );
  MUX2_X1 prince_KeyMUX1_MUXInst_63_U1 ( .A(Key1[64]), .B(Key1[127]), .S(
        prince_KeyMUX1_n8), .Z(prince_selected_Key1_63_) );
  BUF_X1 prince_KeyMUX2_U4 ( .A(prince_n3), .Z(prince_KeyMUX2_n8) );
  BUF_X1 prince_KeyMUX2_U3 ( .A(prince_KeyMUX2_n8), .Z(prince_KeyMUX2_n10) );
  BUF_X1 prince_KeyMUX2_U2 ( .A(prince_n3), .Z(prince_KeyMUX2_n7) );
  BUF_X1 prince_KeyMUX2_U1 ( .A(prince_KeyMUX2_n7), .Z(prince_KeyMUX2_n9) );
  MUX2_X1 prince_KeyMUX2_MUXInst_0_U1 ( .A(prince_k_0_p_share2_0_), .B(
        Key2[64]), .S(prince_KeyMUX2_n7), .Z(prince_selected_Key2_0_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_1_U1 ( .A(Key2[66]), .B(Key2[65]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_1_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_2_U1 ( .A(Key2[67]), .B(Key2[66]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_2_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_3_U1 ( .A(Key2[68]), .B(Key2[67]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_3_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_4_U1 ( .A(Key2[69]), .B(Key2[68]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_4_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_5_U1 ( .A(Key2[70]), .B(Key2[69]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_5_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_6_U1 ( .A(Key2[71]), .B(Key2[70]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_6_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_7_U1 ( .A(Key2[72]), .B(Key2[71]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_7_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_8_U1 ( .A(Key2[73]), .B(Key2[72]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_8_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_9_U1 ( .A(Key2[74]), .B(Key2[73]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_9_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_10_U1 ( .A(Key2[75]), .B(Key2[74]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_10_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_11_U1 ( .A(Key2[76]), .B(Key2[75]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_11_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_12_U1 ( .A(Key2[77]), .B(Key2[76]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_12_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_13_U1 ( .A(Key2[78]), .B(Key2[77]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_13_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_14_U1 ( .A(Key2[79]), .B(Key2[78]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_14_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_15_U1 ( .A(Key2[80]), .B(Key2[79]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_15_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_16_U1 ( .A(Key2[81]), .B(Key2[80]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_16_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_17_U1 ( .A(Key2[82]), .B(Key2[81]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_17_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_18_U1 ( .A(Key2[83]), .B(Key2[82]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_18_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_19_U1 ( .A(Key2[84]), .B(Key2[83]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_19_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_20_U1 ( .A(Key2[85]), .B(Key2[84]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_20_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_21_U1 ( .A(Key2[86]), .B(Key2[85]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_21_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_22_U1 ( .A(Key2[87]), .B(Key2[86]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_22_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_23_U1 ( .A(Key2[88]), .B(Key2[87]), .S(
        prince_KeyMUX2_n7), .Z(prince_selected_Key2_23_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_24_U1 ( .A(Key2[89]), .B(Key2[88]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_24_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_25_U1 ( .A(Key2[90]), .B(Key2[89]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_25_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_26_U1 ( .A(Key2[91]), .B(Key2[90]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_26_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_27_U1 ( .A(Key2[92]), .B(Key2[91]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_27_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_28_U1 ( .A(Key2[93]), .B(Key2[92]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_28_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_29_U1 ( .A(Key2[94]), .B(Key2[93]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_29_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_30_U1 ( .A(Key2[95]), .B(Key2[94]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_30_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_31_U1 ( .A(Key2[96]), .B(Key2[95]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_31_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_32_U1 ( .A(Key2[97]), .B(Key2[96]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_32_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_33_U1 ( .A(Key2[98]), .B(Key2[97]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_33_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_34_U1 ( .A(Key2[99]), .B(Key2[98]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_34_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_35_U1 ( .A(Key2[100]), .B(Key2[99]), .S(
        prince_KeyMUX2_n9), .Z(prince_selected_Key2_35_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_36_U1 ( .A(Key2[101]), .B(Key2[100]), .S(
        prince_KeyMUX2_n10), .Z(prince_selected_Key2_36_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_37_U1 ( .A(Key2[102]), .B(Key2[101]), .S(
        prince_KeyMUX2_n8), .Z(prince_selected_Key2_37_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_38_U1 ( .A(Key2[103]), .B(Key2[102]), .S(
        prince_KeyMUX2_n10), .Z(prince_selected_Key2_38_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_39_U1 ( .A(Key2[104]), .B(Key2[103]), .S(
        prince_KeyMUX2_n8), .Z(prince_selected_Key2_39_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_40_U1 ( .A(Key2[105]), .B(Key2[104]), .S(
        prince_KeyMUX2_n10), .Z(prince_selected_Key2_40_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_41_U1 ( .A(Key2[106]), .B(Key2[105]), .S(
        prince_KeyMUX2_n8), .Z(prince_selected_Key2_41_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_42_U1 ( .A(Key2[107]), .B(Key2[106]), .S(
        prince_KeyMUX2_n8), .Z(prince_selected_Key2_42_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_43_U1 ( .A(Key2[108]), .B(Key2[107]), .S(
        prince_KeyMUX2_n8), .Z(prince_selected_Key2_43_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_44_U1 ( .A(Key2[109]), .B(Key2[108]), .S(
        prince_KeyMUX2_n8), .Z(prince_selected_Key2_44_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_45_U1 ( .A(Key2[110]), .B(Key2[109]), .S(
        prince_KeyMUX2_n8), .Z(prince_selected_Key2_45_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_46_U1 ( .A(Key2[111]), .B(Key2[110]), .S(
        prince_KeyMUX2_n8), .Z(prince_selected_Key2_46_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_47_U1 ( .A(Key2[112]), .B(Key2[111]), .S(
        prince_KeyMUX2_n8), .Z(prince_selected_Key2_47_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_48_U1 ( .A(Key2[113]), .B(Key2[112]), .S(
        prince_KeyMUX2_n10), .Z(prince_selected_Key2_48_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_49_U1 ( .A(Key2[114]), .B(Key2[113]), .S(
        prince_KeyMUX2_n10), .Z(prince_selected_Key2_49_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_50_U1 ( .A(Key2[115]), .B(Key2[114]), .S(
        prince_KeyMUX2_n10), .Z(prince_selected_Key2_50_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_51_U1 ( .A(Key2[116]), .B(Key2[115]), .S(
        prince_KeyMUX2_n10), .Z(prince_selected_Key2_51_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_52_U1 ( .A(Key2[117]), .B(Key2[116]), .S(
        prince_KeyMUX2_n10), .Z(prince_selected_Key2_52_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_53_U1 ( .A(Key2[118]), .B(Key2[117]), .S(
        prince_KeyMUX2_n10), .Z(prince_selected_Key2_53_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_54_U1 ( .A(Key2[119]), .B(Key2[118]), .S(
        prince_KeyMUX2_n10), .Z(prince_selected_Key2_54_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_55_U1 ( .A(Key2[120]), .B(Key2[119]), .S(
        prince_KeyMUX2_n10), .Z(prince_selected_Key2_55_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_56_U1 ( .A(Key2[121]), .B(Key2[120]), .S(
        prince_KeyMUX2_n10), .Z(prince_selected_Key2_56_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_57_U1 ( .A(Key2[122]), .B(Key2[121]), .S(
        prince_KeyMUX2_n10), .Z(prince_selected_Key2_57_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_58_U1 ( .A(Key2[123]), .B(Key2[122]), .S(
        prince_KeyMUX2_n10), .Z(prince_selected_Key2_58_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_59_U1 ( .A(Key2[124]), .B(Key2[123]), .S(
        prince_KeyMUX2_n10), .Z(prince_selected_Key2_59_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_60_U1 ( .A(Key2[125]), .B(Key2[124]), .S(
        prince_KeyMUX2_n8), .Z(prince_selected_Key2_60_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_61_U1 ( .A(Key2[126]), .B(Key2[125]), .S(
        prince_KeyMUX2_n8), .Z(prince_selected_Key2_61_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_62_U1 ( .A(Key2[127]), .B(Key2[126]), .S(
        prince_KeyMUX2_n8), .Z(prince_selected_Key2_62_) );
  MUX2_X1 prince_KeyMUX2_MUXInst_63_U1 ( .A(Key2[64]), .B(Key2[127]), .S(
        prince_KeyMUX2_n8), .Z(prince_selected_Key2_63_) );
  BUF_X1 prince_KeyMUX3_U3 ( .A(prince_n3), .Z(prince_KeyMUX3_n7) );
  BUF_X1 prince_KeyMUX3_U2 ( .A(prince_KeyMUX3_n7), .Z(prince_KeyMUX3_n9) );
  BUF_X1 prince_KeyMUX3_U1 ( .A(prince_n3), .Z(prince_KeyMUX3_n8) );
  MUX2_X1 prince_KeyMUX3_MUXInst_0_U1 ( .A(prince_k_0_p_share3_0_), .B(
        Key3[64]), .S(prince_n3), .Z(prince_selected_Key3_0_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_1_U1 ( .A(Key3[66]), .B(Key3[65]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_1_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_2_U1 ( .A(Key3[67]), .B(Key3[66]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_2_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_3_U1 ( .A(Key3[68]), .B(Key3[67]), .S(
        prince_n3), .Z(prince_selected_Key3_3_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_4_U1 ( .A(Key3[69]), .B(Key3[68]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_4_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_5_U1 ( .A(Key3[70]), .B(Key3[69]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_5_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_6_U1 ( .A(Key3[71]), .B(Key3[70]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_6_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_7_U1 ( .A(Key3[72]), .B(Key3[71]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_7_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_8_U1 ( .A(Key3[73]), .B(Key3[72]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_8_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_9_U1 ( .A(Key3[74]), .B(Key3[73]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_9_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_10_U1 ( .A(Key3[75]), .B(Key3[74]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_10_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_11_U1 ( .A(Key3[76]), .B(Key3[75]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_11_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_12_U1 ( .A(Key3[77]), .B(Key3[76]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_12_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_13_U1 ( .A(Key3[78]), .B(Key3[77]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_13_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_14_U1 ( .A(Key3[79]), .B(Key3[78]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_14_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_15_U1 ( .A(Key3[80]), .B(Key3[79]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_15_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_16_U1 ( .A(Key3[81]), .B(Key3[80]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_16_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_17_U1 ( .A(Key3[82]), .B(Key3[81]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_17_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_18_U1 ( .A(Key3[83]), .B(Key3[82]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_18_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_19_U1 ( .A(Key3[84]), .B(Key3[83]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_19_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_20_U1 ( .A(Key3[85]), .B(Key3[84]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_20_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_21_U1 ( .A(Key3[86]), .B(Key3[85]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_21_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_22_U1 ( .A(Key3[87]), .B(Key3[86]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_22_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_23_U1 ( .A(Key3[88]), .B(Key3[87]), .S(
        prince_KeyMUX3_n7), .Z(prince_selected_Key3_23_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_24_U1 ( .A(Key3[89]), .B(Key3[88]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_24_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_25_U1 ( .A(Key3[90]), .B(Key3[89]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_25_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_26_U1 ( .A(Key3[91]), .B(Key3[90]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_26_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_27_U1 ( .A(Key3[92]), .B(Key3[91]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_27_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_28_U1 ( .A(Key3[93]), .B(Key3[92]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_28_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_29_U1 ( .A(Key3[94]), .B(Key3[93]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_29_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_30_U1 ( .A(Key3[95]), .B(Key3[94]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_30_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_31_U1 ( .A(Key3[96]), .B(Key3[95]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_31_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_32_U1 ( .A(Key3[97]), .B(Key3[96]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_32_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_33_U1 ( .A(Key3[98]), .B(Key3[97]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_33_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_34_U1 ( .A(Key3[99]), .B(Key3[98]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_34_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_35_U1 ( .A(Key3[100]), .B(Key3[99]), .S(
        prince_KeyMUX3_n9), .Z(prince_selected_Key3_35_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_36_U1 ( .A(Key3[101]), .B(Key3[100]), .S(
        prince_KeyMUX3_n8), .Z(prince_selected_Key3_36_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_37_U1 ( .A(Key3[102]), .B(Key3[101]), .S(
        prince_n3), .Z(prince_selected_Key3_37_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_38_U1 ( .A(Key3[103]), .B(Key3[102]), .S(
        prince_KeyMUX3_n8), .Z(prince_selected_Key3_38_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_39_U1 ( .A(Key3[104]), .B(Key3[103]), .S(
        prince_n3), .Z(prince_selected_Key3_39_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_40_U1 ( .A(Key3[105]), .B(Key3[104]), .S(
        prince_KeyMUX3_n8), .Z(prince_selected_Key3_40_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_41_U1 ( .A(Key3[106]), .B(Key3[105]), .S(
        prince_n3), .Z(prince_selected_Key3_41_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_42_U1 ( .A(Key3[107]), .B(Key3[106]), .S(
        prince_KeyMUX3_n8), .Z(prince_selected_Key3_42_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_43_U1 ( .A(Key3[108]), .B(Key3[107]), .S(
        prince_n3), .Z(prince_selected_Key3_43_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_44_U1 ( .A(Key3[109]), .B(Key3[108]), .S(
        prince_KeyMUX3_n8), .Z(prince_selected_Key3_44_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_45_U1 ( .A(Key3[110]), .B(Key3[109]), .S(
        prince_n3), .Z(prince_selected_Key3_45_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_46_U1 ( .A(Key3[111]), .B(Key3[110]), .S(
        prince_KeyMUX3_n8), .Z(prince_selected_Key3_46_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_47_U1 ( .A(Key3[112]), .B(Key3[111]), .S(
        prince_KeyMUX3_n8), .Z(prince_selected_Key3_47_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_48_U1 ( .A(Key3[113]), .B(Key3[112]), .S(
        prince_KeyMUX3_n8), .Z(prince_selected_Key3_48_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_49_U1 ( .A(Key3[114]), .B(Key3[113]), .S(
        prince_n3), .Z(prince_selected_Key3_49_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_50_U1 ( .A(Key3[115]), .B(Key3[114]), .S(
        prince_KeyMUX3_n8), .Z(prince_selected_Key3_50_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_51_U1 ( .A(Key3[116]), .B(Key3[115]), .S(
        prince_n3), .Z(prince_selected_Key3_51_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_52_U1 ( .A(Key3[117]), .B(Key3[116]), .S(
        prince_KeyMUX3_n8), .Z(prince_selected_Key3_52_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_53_U1 ( .A(Key3[118]), .B(Key3[117]), .S(
        prince_n3), .Z(prince_selected_Key3_53_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_54_U1 ( .A(Key3[119]), .B(Key3[118]), .S(
        prince_KeyMUX3_n8), .Z(prince_selected_Key3_54_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_55_U1 ( .A(Key3[120]), .B(Key3[119]), .S(
        prince_n3), .Z(prince_selected_Key3_55_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_56_U1 ( .A(Key3[121]), .B(Key3[120]), .S(
        prince_KeyMUX3_n8), .Z(prince_selected_Key3_56_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_57_U1 ( .A(Key3[122]), .B(Key3[121]), .S(
        prince_n3), .Z(prince_selected_Key3_57_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_58_U1 ( .A(Key3[123]), .B(Key3[122]), .S(
        prince_KeyMUX3_n8), .Z(prince_selected_Key3_58_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_59_U1 ( .A(Key3[124]), .B(Key3[123]), .S(
        prince_KeyMUX3_n8), .Z(prince_selected_Key3_59_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_60_U1 ( .A(Key3[125]), .B(Key3[124]), .S(
        prince_n3), .Z(prince_selected_Key3_60_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_61_U1 ( .A(Key3[126]), .B(Key3[125]), .S(
        prince_KeyMUX3_n8), .Z(prince_selected_Key3_61_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_62_U1 ( .A(Key3[127]), .B(Key3[126]), .S(
        prince_n3), .Z(prince_selected_Key3_62_) );
  MUX2_X1 prince_KeyMUX3_MUXInst_63_U1 ( .A(Key3[64]), .B(Key3[127]), .S(
        prince_KeyMUX3_n8), .Z(prince_selected_Key3_63_) );
  XNOR2_X1 prince_AddKey1_XORInst_0_0_U2 ( .A(prince_AddKey1_XORInst_0_0_n3), 
        .B(prince_selected_Key1_0_), .ZN(prince_SR_Inv_Result_s1[16]) );
  XNOR2_X1 prince_AddKey1_XORInst_0_0_U1 ( .A(1'b0), .B(input_s1[0]), .ZN(
        prince_AddKey1_XORInst_0_0_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_0_1_U2 ( .A(prince_AddKey1_XORInst_0_1_n3), 
        .B(prince_selected_Key1_1_), .ZN(prince_SR_Inv_Result_s1[17]) );
  XNOR2_X1 prince_AddKey1_XORInst_0_1_U1 ( .A(1'b0), .B(input_s1[1]), .ZN(
        prince_AddKey1_XORInst_0_1_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_0_2_U2 ( .A(prince_AddKey1_XORInst_0_2_n3), 
        .B(prince_selected_Key1_2_), .ZN(prince_SR_Inv_Result_s1[18]) );
  XNOR2_X1 prince_AddKey1_XORInst_0_2_U1 ( .A(1'b0), .B(input_s1[2]), .ZN(
        prince_AddKey1_XORInst_0_2_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_0_3_U2 ( .A(prince_AddKey1_XORInst_0_3_n3), 
        .B(prince_selected_Key1_3_), .ZN(prince_SR_Inv_Result_s1[19]) );
  XNOR2_X1 prince_AddKey1_XORInst_0_3_U1 ( .A(1'b0), .B(input_s1[3]), .ZN(
        prince_AddKey1_XORInst_0_3_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_1_0_U2 ( .A(prince_AddKey1_XORInst_1_0_n3), 
        .B(prince_selected_Key1_4_), .ZN(prince_SR_Inv_Result_s1[36]) );
  XNOR2_X1 prince_AddKey1_XORInst_1_0_U1 ( .A(1'b0), .B(input_s1[4]), .ZN(
        prince_AddKey1_XORInst_1_0_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_1_1_U2 ( .A(prince_AddKey1_XORInst_1_1_n3), 
        .B(prince_selected_Key1_5_), .ZN(prince_SR_Inv_Result_s1[37]) );
  XNOR2_X1 prince_AddKey1_XORInst_1_1_U1 ( .A(1'b0), .B(input_s1[5]), .ZN(
        prince_AddKey1_XORInst_1_1_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_1_2_U2 ( .A(prince_AddKey1_XORInst_1_2_n3), 
        .B(prince_selected_Key1_6_), .ZN(prince_SR_Inv_Result_s1[38]) );
  XNOR2_X1 prince_AddKey1_XORInst_1_2_U1 ( .A(1'b0), .B(input_s1[6]), .ZN(
        prince_AddKey1_XORInst_1_2_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_1_3_U2 ( .A(prince_AddKey1_XORInst_1_3_n3), 
        .B(prince_selected_Key1_7_), .ZN(prince_SR_Inv_Result_s1[39]) );
  XNOR2_X1 prince_AddKey1_XORInst_1_3_U1 ( .A(1'b0), .B(input_s1[7]), .ZN(
        prince_AddKey1_XORInst_1_3_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_2_0_U2 ( .A(prince_AddKey1_XORInst_2_0_n3), 
        .B(prince_selected_Key1_8_), .ZN(prince_SR_Inv_Result_s1[56]) );
  XNOR2_X1 prince_AddKey1_XORInst_2_0_U1 ( .A(1'b0), .B(input_s1[8]), .ZN(
        prince_AddKey1_XORInst_2_0_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_2_1_U2 ( .A(prince_AddKey1_XORInst_2_1_n3), 
        .B(prince_selected_Key1_9_), .ZN(prince_SR_Inv_Result_s1[57]) );
  XNOR2_X1 prince_AddKey1_XORInst_2_1_U1 ( .A(1'b0), .B(input_s1[9]), .ZN(
        prince_AddKey1_XORInst_2_1_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_2_2_U2 ( .A(prince_AddKey1_XORInst_2_2_n3), 
        .B(prince_selected_Key1_10_), .ZN(prince_SR_Inv_Result_s1[58]) );
  XNOR2_X1 prince_AddKey1_XORInst_2_2_U1 ( .A(1'b0), .B(input_s1[10]), .ZN(
        prince_AddKey1_XORInst_2_2_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_2_3_U2 ( .A(prince_AddKey1_XORInst_2_3_n3), 
        .B(prince_selected_Key1_11_), .ZN(prince_SR_Inv_Result_s1[59]) );
  XNOR2_X1 prince_AddKey1_XORInst_2_3_U1 ( .A(1'b0), .B(input_s1[11]), .ZN(
        prince_AddKey1_XORInst_2_3_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_3_0_U2 ( .A(prince_AddKey1_XORInst_3_0_n3), 
        .B(prince_selected_Key1_12_), .ZN(prince_SR_Inv_Result_s1[12]) );
  XNOR2_X1 prince_AddKey1_XORInst_3_0_U1 ( .A(1'b0), .B(input_s1[12]), .ZN(
        prince_AddKey1_XORInst_3_0_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_3_1_U2 ( .A(prince_AddKey1_XORInst_3_1_n3), 
        .B(prince_selected_Key1_13_), .ZN(prince_SR_Inv_Result_s1[13]) );
  XNOR2_X1 prince_AddKey1_XORInst_3_1_U1 ( .A(1'b0), .B(input_s1[13]), .ZN(
        prince_AddKey1_XORInst_3_1_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_3_2_U2 ( .A(prince_AddKey1_XORInst_3_2_n3), 
        .B(prince_selected_Key1_14_), .ZN(prince_SR_Inv_Result_s1[14]) );
  XNOR2_X1 prince_AddKey1_XORInst_3_2_U1 ( .A(1'b0), .B(input_s1[14]), .ZN(
        prince_AddKey1_XORInst_3_2_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_3_3_U2 ( .A(prince_AddKey1_XORInst_3_3_n3), 
        .B(prince_selected_Key1_15_), .ZN(prince_SR_Inv_Result_s1[15]) );
  XNOR2_X1 prince_AddKey1_XORInst_3_3_U1 ( .A(1'b0), .B(input_s1[15]), .ZN(
        prince_AddKey1_XORInst_3_3_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_4_0_U2 ( .A(prince_AddKey1_XORInst_4_0_n3), 
        .B(prince_selected_Key1_16_), .ZN(prince_SR_Inv_Result_s1[32]) );
  XNOR2_X1 prince_AddKey1_XORInst_4_0_U1 ( .A(1'b0), .B(input_s1[16]), .ZN(
        prince_AddKey1_XORInst_4_0_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_4_1_U2 ( .A(prince_AddKey1_XORInst_4_1_n3), 
        .B(prince_selected_Key1_17_), .ZN(prince_SR_Inv_Result_s1[33]) );
  XNOR2_X1 prince_AddKey1_XORInst_4_1_U1 ( .A(1'b0), .B(input_s1[17]), .ZN(
        prince_AddKey1_XORInst_4_1_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_4_2_U2 ( .A(prince_AddKey1_XORInst_4_2_n3), 
        .B(prince_selected_Key1_18_), .ZN(prince_SR_Inv_Result_s1[34]) );
  XNOR2_X1 prince_AddKey1_XORInst_4_2_U1 ( .A(1'b0), .B(input_s1[18]), .ZN(
        prince_AddKey1_XORInst_4_2_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_4_3_U2 ( .A(prince_AddKey1_XORInst_4_3_n3), 
        .B(prince_selected_Key1_19_), .ZN(prince_SR_Inv_Result_s1[35]) );
  XNOR2_X1 prince_AddKey1_XORInst_4_3_U1 ( .A(1'b0), .B(input_s1[19]), .ZN(
        prince_AddKey1_XORInst_4_3_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_5_0_U2 ( .A(prince_AddKey1_XORInst_5_0_n3), 
        .B(prince_selected_Key1_20_), .ZN(prince_SR_Inv_Result_s1[52]) );
  XNOR2_X1 prince_AddKey1_XORInst_5_0_U1 ( .A(1'b0), .B(input_s1[20]), .ZN(
        prince_AddKey1_XORInst_5_0_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_5_1_U2 ( .A(prince_AddKey1_XORInst_5_1_n3), 
        .B(prince_selected_Key1_21_), .ZN(prince_SR_Inv_Result_s1[53]) );
  XNOR2_X1 prince_AddKey1_XORInst_5_1_U1 ( .A(1'b0), .B(input_s1[21]), .ZN(
        prince_AddKey1_XORInst_5_1_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_5_2_U2 ( .A(prince_AddKey1_XORInst_5_2_n3), 
        .B(prince_selected_Key1_22_), .ZN(prince_SR_Inv_Result_s1[54]) );
  XNOR2_X1 prince_AddKey1_XORInst_5_2_U1 ( .A(1'b0), .B(input_s1[22]), .ZN(
        prince_AddKey1_XORInst_5_2_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_5_3_U2 ( .A(prince_AddKey1_XORInst_5_3_n3), 
        .B(prince_selected_Key1_23_), .ZN(prince_SR_Inv_Result_s1[55]) );
  XNOR2_X1 prince_AddKey1_XORInst_5_3_U1 ( .A(1'b0), .B(input_s1[23]), .ZN(
        prince_AddKey1_XORInst_5_3_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_6_0_U2 ( .A(prince_AddKey1_XORInst_6_0_n3), 
        .B(prince_selected_Key1_24_), .ZN(prince_SR_Inv_Result_s1[8]) );
  XNOR2_X1 prince_AddKey1_XORInst_6_0_U1 ( .A(1'b0), .B(input_s1[24]), .ZN(
        prince_AddKey1_XORInst_6_0_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_6_1_U2 ( .A(prince_AddKey1_XORInst_6_1_n3), 
        .B(prince_selected_Key1_25_), .ZN(prince_SR_Inv_Result_s1[9]) );
  XNOR2_X1 prince_AddKey1_XORInst_6_1_U1 ( .A(1'b0), .B(input_s1[25]), .ZN(
        prince_AddKey1_XORInst_6_1_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_6_2_U2 ( .A(prince_AddKey1_XORInst_6_2_n3), 
        .B(prince_selected_Key1_26_), .ZN(prince_SR_Inv_Result_s1[10]) );
  XNOR2_X1 prince_AddKey1_XORInst_6_2_U1 ( .A(1'b0), .B(input_s1[26]), .ZN(
        prince_AddKey1_XORInst_6_2_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_6_3_U2 ( .A(prince_AddKey1_XORInst_6_3_n3), 
        .B(prince_selected_Key1_27_), .ZN(prince_SR_Inv_Result_s1[11]) );
  XNOR2_X1 prince_AddKey1_XORInst_6_3_U1 ( .A(1'b0), .B(input_s1[27]), .ZN(
        prince_AddKey1_XORInst_6_3_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_7_0_U2 ( .A(prince_AddKey1_XORInst_7_0_n3), 
        .B(prince_selected_Key1_28_), .ZN(prince_SR_Inv_Result_s1[28]) );
  XNOR2_X1 prince_AddKey1_XORInst_7_0_U1 ( .A(1'b0), .B(input_s1[28]), .ZN(
        prince_AddKey1_XORInst_7_0_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_7_1_U2 ( .A(prince_AddKey1_XORInst_7_1_n3), 
        .B(prince_selected_Key1_29_), .ZN(prince_SR_Inv_Result_s1[29]) );
  XNOR2_X1 prince_AddKey1_XORInst_7_1_U1 ( .A(1'b0), .B(input_s1[29]), .ZN(
        prince_AddKey1_XORInst_7_1_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_7_2_U2 ( .A(prince_AddKey1_XORInst_7_2_n3), 
        .B(prince_selected_Key1_30_), .ZN(prince_SR_Inv_Result_s1[30]) );
  XNOR2_X1 prince_AddKey1_XORInst_7_2_U1 ( .A(1'b0), .B(input_s1[30]), .ZN(
        prince_AddKey1_XORInst_7_2_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_7_3_U2 ( .A(prince_AddKey1_XORInst_7_3_n3), 
        .B(prince_selected_Key1_31_), .ZN(prince_SR_Inv_Result_s1[31]) );
  XNOR2_X1 prince_AddKey1_XORInst_7_3_U1 ( .A(1'b0), .B(input_s1[31]), .ZN(
        prince_AddKey1_XORInst_7_3_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_8_0_U2 ( .A(prince_AddKey1_XORInst_8_0_n3), 
        .B(prince_selected_Key1_32_), .ZN(prince_SR_Inv_Result_s1[48]) );
  XNOR2_X1 prince_AddKey1_XORInst_8_0_U1 ( .A(1'b0), .B(input_s1[32]), .ZN(
        prince_AddKey1_XORInst_8_0_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_8_1_U2 ( .A(prince_AddKey1_XORInst_8_1_n3), 
        .B(prince_selected_Key1_33_), .ZN(prince_SR_Inv_Result_s1[49]) );
  XNOR2_X1 prince_AddKey1_XORInst_8_1_U1 ( .A(1'b0), .B(input_s1[33]), .ZN(
        prince_AddKey1_XORInst_8_1_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_8_2_U2 ( .A(prince_AddKey1_XORInst_8_2_n3), 
        .B(prince_selected_Key1_34_), .ZN(prince_SR_Inv_Result_s1[50]) );
  XNOR2_X1 prince_AddKey1_XORInst_8_2_U1 ( .A(1'b0), .B(input_s1[34]), .ZN(
        prince_AddKey1_XORInst_8_2_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_8_3_U2 ( .A(prince_AddKey1_XORInst_8_3_n3), 
        .B(prince_selected_Key1_35_), .ZN(prince_SR_Inv_Result_s1[51]) );
  XNOR2_X1 prince_AddKey1_XORInst_8_3_U1 ( .A(1'b0), .B(input_s1[35]), .ZN(
        prince_AddKey1_XORInst_8_3_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_9_0_U2 ( .A(prince_AddKey1_XORInst_9_0_n3), 
        .B(prince_selected_Key1_36_), .ZN(prince_SR_Inv_Result_s1[4]) );
  XNOR2_X1 prince_AddKey1_XORInst_9_0_U1 ( .A(1'b0), .B(input_s1[36]), .ZN(
        prince_AddKey1_XORInst_9_0_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_9_1_U2 ( .A(prince_AddKey1_XORInst_9_1_n3), 
        .B(prince_selected_Key1_37_), .ZN(prince_SR_Inv_Result_s1[5]) );
  XNOR2_X1 prince_AddKey1_XORInst_9_1_U1 ( .A(1'b0), .B(input_s1[37]), .ZN(
        prince_AddKey1_XORInst_9_1_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_9_2_U2 ( .A(prince_AddKey1_XORInst_9_2_n3), 
        .B(prince_selected_Key1_38_), .ZN(prince_SR_Inv_Result_s1[6]) );
  XNOR2_X1 prince_AddKey1_XORInst_9_2_U1 ( .A(1'b0), .B(input_s1[38]), .ZN(
        prince_AddKey1_XORInst_9_2_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_9_3_U2 ( .A(prince_AddKey1_XORInst_9_3_n3), 
        .B(prince_selected_Key1_39_), .ZN(prince_SR_Inv_Result_s1[7]) );
  XNOR2_X1 prince_AddKey1_XORInst_9_3_U1 ( .A(1'b0), .B(input_s1[39]), .ZN(
        prince_AddKey1_XORInst_9_3_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_10_0_U2 ( .A(prince_AddKey1_XORInst_10_0_n3), 
        .B(prince_selected_Key1_40_), .ZN(prince_SR_Inv_Result_s1[24]) );
  XNOR2_X1 prince_AddKey1_XORInst_10_0_U1 ( .A(1'b0), .B(input_s1[40]), .ZN(
        prince_AddKey1_XORInst_10_0_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_10_1_U2 ( .A(prince_AddKey1_XORInst_10_1_n3), 
        .B(prince_selected_Key1_41_), .ZN(prince_SR_Inv_Result_s1[25]) );
  XNOR2_X1 prince_AddKey1_XORInst_10_1_U1 ( .A(1'b0), .B(input_s1[41]), .ZN(
        prince_AddKey1_XORInst_10_1_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_10_2_U2 ( .A(prince_AddKey1_XORInst_10_2_n3), 
        .B(prince_selected_Key1_42_), .ZN(prince_SR_Inv_Result_s1[26]) );
  XNOR2_X1 prince_AddKey1_XORInst_10_2_U1 ( .A(1'b0), .B(input_s1[42]), .ZN(
        prince_AddKey1_XORInst_10_2_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_10_3_U2 ( .A(prince_AddKey1_XORInst_10_3_n3), 
        .B(prince_selected_Key1_43_), .ZN(prince_SR_Inv_Result_s1[27]) );
  XNOR2_X1 prince_AddKey1_XORInst_10_3_U1 ( .A(1'b0), .B(input_s1[43]), .ZN(
        prince_AddKey1_XORInst_10_3_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_11_0_U2 ( .A(prince_AddKey1_XORInst_11_0_n3), 
        .B(prince_selected_Key1_44_), .ZN(prince_SR_Inv_Result_s1[44]) );
  XNOR2_X1 prince_AddKey1_XORInst_11_0_U1 ( .A(1'b0), .B(input_s1[44]), .ZN(
        prince_AddKey1_XORInst_11_0_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_11_1_U2 ( .A(prince_AddKey1_XORInst_11_1_n3), 
        .B(prince_selected_Key1_45_), .ZN(prince_SR_Inv_Result_s1[45]) );
  XNOR2_X1 prince_AddKey1_XORInst_11_1_U1 ( .A(1'b0), .B(input_s1[45]), .ZN(
        prince_AddKey1_XORInst_11_1_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_11_2_U2 ( .A(prince_AddKey1_XORInst_11_2_n3), 
        .B(prince_selected_Key1_46_), .ZN(prince_SR_Inv_Result_s1[46]) );
  XNOR2_X1 prince_AddKey1_XORInst_11_2_U1 ( .A(1'b0), .B(input_s1[46]), .ZN(
        prince_AddKey1_XORInst_11_2_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_11_3_U2 ( .A(prince_AddKey1_XORInst_11_3_n3), 
        .B(prince_selected_Key1_47_), .ZN(prince_SR_Inv_Result_s1[47]) );
  XNOR2_X1 prince_AddKey1_XORInst_11_3_U1 ( .A(1'b0), .B(input_s1[47]), .ZN(
        prince_AddKey1_XORInst_11_3_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_12_0_U2 ( .A(prince_AddKey1_XORInst_12_0_n3), 
        .B(prince_selected_Key1_48_), .ZN(prince_SR_Inv_Result_s1[0]) );
  XNOR2_X1 prince_AddKey1_XORInst_12_0_U1 ( .A(1'b0), .B(input_s1[48]), .ZN(
        prince_AddKey1_XORInst_12_0_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_12_1_U2 ( .A(prince_AddKey1_XORInst_12_1_n3), 
        .B(prince_selected_Key1_49_), .ZN(prince_SR_Inv_Result_s1[1]) );
  XNOR2_X1 prince_AddKey1_XORInst_12_1_U1 ( .A(1'b0), .B(input_s1[49]), .ZN(
        prince_AddKey1_XORInst_12_1_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_12_2_U2 ( .A(prince_AddKey1_XORInst_12_2_n3), 
        .B(prince_selected_Key1_50_), .ZN(prince_SR_Inv_Result_s1[2]) );
  XNOR2_X1 prince_AddKey1_XORInst_12_2_U1 ( .A(1'b0), .B(input_s1[50]), .ZN(
        prince_AddKey1_XORInst_12_2_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_12_3_U2 ( .A(prince_AddKey1_XORInst_12_3_n3), 
        .B(prince_selected_Key1_51_), .ZN(prince_SR_Inv_Result_s1[3]) );
  XNOR2_X1 prince_AddKey1_XORInst_12_3_U1 ( .A(1'b0), .B(input_s1[51]), .ZN(
        prince_AddKey1_XORInst_12_3_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_13_0_U2 ( .A(prince_AddKey1_XORInst_13_0_n3), 
        .B(prince_selected_Key1_52_), .ZN(prince_SR_Inv_Result_s1[20]) );
  XNOR2_X1 prince_AddKey1_XORInst_13_0_U1 ( .A(1'b0), .B(input_s1[52]), .ZN(
        prince_AddKey1_XORInst_13_0_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_13_1_U2 ( .A(prince_AddKey1_XORInst_13_1_n3), 
        .B(prince_selected_Key1_53_), .ZN(prince_SR_Inv_Result_s1[21]) );
  XNOR2_X1 prince_AddKey1_XORInst_13_1_U1 ( .A(1'b0), .B(input_s1[53]), .ZN(
        prince_AddKey1_XORInst_13_1_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_13_2_U2 ( .A(prince_AddKey1_XORInst_13_2_n3), 
        .B(prince_selected_Key1_54_), .ZN(prince_SR_Inv_Result_s1[22]) );
  XNOR2_X1 prince_AddKey1_XORInst_13_2_U1 ( .A(1'b0), .B(input_s1[54]), .ZN(
        prince_AddKey1_XORInst_13_2_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_13_3_U2 ( .A(prince_AddKey1_XORInst_13_3_n3), 
        .B(prince_selected_Key1_55_), .ZN(prince_SR_Inv_Result_s1[23]) );
  XNOR2_X1 prince_AddKey1_XORInst_13_3_U1 ( .A(1'b0), .B(input_s1[55]), .ZN(
        prince_AddKey1_XORInst_13_3_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_14_0_U2 ( .A(prince_AddKey1_XORInst_14_0_n3), 
        .B(prince_selected_Key1_56_), .ZN(prince_SR_Inv_Result_s1[40]) );
  XNOR2_X1 prince_AddKey1_XORInst_14_0_U1 ( .A(1'b0), .B(input_s1[56]), .ZN(
        prince_AddKey1_XORInst_14_0_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_14_1_U2 ( .A(prince_AddKey1_XORInst_14_1_n3), 
        .B(prince_selected_Key1_57_), .ZN(prince_SR_Inv_Result_s1[41]) );
  XNOR2_X1 prince_AddKey1_XORInst_14_1_U1 ( .A(1'b0), .B(input_s1[57]), .ZN(
        prince_AddKey1_XORInst_14_1_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_14_2_U2 ( .A(prince_AddKey1_XORInst_14_2_n3), 
        .B(prince_selected_Key1_58_), .ZN(prince_SR_Inv_Result_s1[42]) );
  XNOR2_X1 prince_AddKey1_XORInst_14_2_U1 ( .A(1'b0), .B(input_s1[58]), .ZN(
        prince_AddKey1_XORInst_14_2_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_14_3_U2 ( .A(prince_AddKey1_XORInst_14_3_n3), 
        .B(prince_selected_Key1_59_), .ZN(prince_SR_Inv_Result_s1[43]) );
  XNOR2_X1 prince_AddKey1_XORInst_14_3_U1 ( .A(1'b0), .B(input_s1[59]), .ZN(
        prince_AddKey1_XORInst_14_3_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_15_0_U2 ( .A(prince_AddKey1_XORInst_15_0_n3), 
        .B(prince_selected_Key1_60_), .ZN(prince_SR_Inv_Result_s1[60]) );
  XNOR2_X1 prince_AddKey1_XORInst_15_0_U1 ( .A(1'b0), .B(input_s1[60]), .ZN(
        prince_AddKey1_XORInst_15_0_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_15_1_U2 ( .A(prince_AddKey1_XORInst_15_1_n3), 
        .B(prince_selected_Key1_61_), .ZN(prince_SR_Inv_Result_s1[61]) );
  XNOR2_X1 prince_AddKey1_XORInst_15_1_U1 ( .A(1'b0), .B(input_s1[61]), .ZN(
        prince_AddKey1_XORInst_15_1_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_15_2_U2 ( .A(prince_AddKey1_XORInst_15_2_n3), 
        .B(prince_selected_Key1_62_), .ZN(prince_SR_Inv_Result_s1[62]) );
  XNOR2_X1 prince_AddKey1_XORInst_15_2_U1 ( .A(1'b0), .B(input_s1[62]), .ZN(
        prince_AddKey1_XORInst_15_2_n3) );
  XNOR2_X1 prince_AddKey1_XORInst_15_3_U2 ( .A(prince_AddKey1_XORInst_15_3_n3), 
        .B(prince_selected_Key1_63_), .ZN(prince_SR_Inv_Result_s1[63]) );
  XNOR2_X1 prince_AddKey1_XORInst_15_3_U1 ( .A(1'b0), .B(input_s1[63]), .ZN(
        prince_AddKey1_XORInst_15_3_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_0_0_U2 ( .A(prince_AddKey2_XORInst_0_0_n3), 
        .B(prince_selected_Key2_0_), .ZN(prince_SR_Inv_Result_s2[16]) );
  XNOR2_X1 prince_AddKey2_XORInst_0_0_U1 ( .A(1'b0), .B(input_s2[0]), .ZN(
        prince_AddKey2_XORInst_0_0_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_0_1_U2 ( .A(prince_AddKey2_XORInst_0_1_n3), 
        .B(prince_selected_Key2_1_), .ZN(prince_SR_Inv_Result_s2[17]) );
  XNOR2_X1 prince_AddKey2_XORInst_0_1_U1 ( .A(1'b0), .B(input_s2[1]), .ZN(
        prince_AddKey2_XORInst_0_1_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_0_2_U2 ( .A(prince_AddKey2_XORInst_0_2_n3), 
        .B(prince_selected_Key2_2_), .ZN(prince_SR_Inv_Result_s2[18]) );
  XNOR2_X1 prince_AddKey2_XORInst_0_2_U1 ( .A(1'b0), .B(input_s2[2]), .ZN(
        prince_AddKey2_XORInst_0_2_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_0_3_U2 ( .A(prince_AddKey2_XORInst_0_3_n3), 
        .B(prince_selected_Key2_3_), .ZN(prince_SR_Inv_Result_s2[19]) );
  XNOR2_X1 prince_AddKey2_XORInst_0_3_U1 ( .A(1'b0), .B(input_s2[3]), .ZN(
        prince_AddKey2_XORInst_0_3_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_1_0_U2 ( .A(prince_AddKey2_XORInst_1_0_n3), 
        .B(prince_selected_Key2_4_), .ZN(prince_SR_Inv_Result_s2[36]) );
  XNOR2_X1 prince_AddKey2_XORInst_1_0_U1 ( .A(1'b0), .B(input_s2[4]), .ZN(
        prince_AddKey2_XORInst_1_0_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_1_1_U2 ( .A(prince_AddKey2_XORInst_1_1_n3), 
        .B(prince_selected_Key2_5_), .ZN(prince_SR_Inv_Result_s2[37]) );
  XNOR2_X1 prince_AddKey2_XORInst_1_1_U1 ( .A(1'b0), .B(input_s2[5]), .ZN(
        prince_AddKey2_XORInst_1_1_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_1_2_U2 ( .A(prince_AddKey2_XORInst_1_2_n3), 
        .B(prince_selected_Key2_6_), .ZN(prince_SR_Inv_Result_s2[38]) );
  XNOR2_X1 prince_AddKey2_XORInst_1_2_U1 ( .A(1'b0), .B(input_s2[6]), .ZN(
        prince_AddKey2_XORInst_1_2_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_1_3_U2 ( .A(prince_AddKey2_XORInst_1_3_n3), 
        .B(prince_selected_Key2_7_), .ZN(prince_SR_Inv_Result_s2[39]) );
  XNOR2_X1 prince_AddKey2_XORInst_1_3_U1 ( .A(1'b0), .B(input_s2[7]), .ZN(
        prince_AddKey2_XORInst_1_3_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_2_0_U2 ( .A(prince_AddKey2_XORInst_2_0_n3), 
        .B(prince_selected_Key2_8_), .ZN(prince_SR_Inv_Result_s2[56]) );
  XNOR2_X1 prince_AddKey2_XORInst_2_0_U1 ( .A(1'b0), .B(input_s2[8]), .ZN(
        prince_AddKey2_XORInst_2_0_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_2_1_U2 ( .A(prince_AddKey2_XORInst_2_1_n3), 
        .B(prince_selected_Key2_9_), .ZN(prince_SR_Inv_Result_s2[57]) );
  XNOR2_X1 prince_AddKey2_XORInst_2_1_U1 ( .A(1'b0), .B(input_s2[9]), .ZN(
        prince_AddKey2_XORInst_2_1_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_2_2_U2 ( .A(prince_AddKey2_XORInst_2_2_n3), 
        .B(prince_selected_Key2_10_), .ZN(prince_SR_Inv_Result_s2[58]) );
  XNOR2_X1 prince_AddKey2_XORInst_2_2_U1 ( .A(1'b0), .B(input_s2[10]), .ZN(
        prince_AddKey2_XORInst_2_2_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_2_3_U2 ( .A(prince_AddKey2_XORInst_2_3_n3), 
        .B(prince_selected_Key2_11_), .ZN(prince_SR_Inv_Result_s2[59]) );
  XNOR2_X1 prince_AddKey2_XORInst_2_3_U1 ( .A(1'b0), .B(input_s2[11]), .ZN(
        prince_AddKey2_XORInst_2_3_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_3_0_U2 ( .A(prince_AddKey2_XORInst_3_0_n3), 
        .B(prince_selected_Key2_12_), .ZN(prince_SR_Inv_Result_s2[12]) );
  XNOR2_X1 prince_AddKey2_XORInst_3_0_U1 ( .A(1'b0), .B(input_s2[12]), .ZN(
        prince_AddKey2_XORInst_3_0_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_3_1_U2 ( .A(prince_AddKey2_XORInst_3_1_n3), 
        .B(prince_selected_Key2_13_), .ZN(prince_SR_Inv_Result_s2[13]) );
  XNOR2_X1 prince_AddKey2_XORInst_3_1_U1 ( .A(1'b0), .B(input_s2[13]), .ZN(
        prince_AddKey2_XORInst_3_1_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_3_2_U2 ( .A(prince_AddKey2_XORInst_3_2_n3), 
        .B(prince_selected_Key2_14_), .ZN(prince_SR_Inv_Result_s2[14]) );
  XNOR2_X1 prince_AddKey2_XORInst_3_2_U1 ( .A(1'b0), .B(input_s2[14]), .ZN(
        prince_AddKey2_XORInst_3_2_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_3_3_U2 ( .A(prince_AddKey2_XORInst_3_3_n3), 
        .B(prince_selected_Key2_15_), .ZN(prince_SR_Inv_Result_s2[15]) );
  XNOR2_X1 prince_AddKey2_XORInst_3_3_U1 ( .A(1'b0), .B(input_s2[15]), .ZN(
        prince_AddKey2_XORInst_3_3_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_4_0_U2 ( .A(prince_AddKey2_XORInst_4_0_n3), 
        .B(prince_selected_Key2_16_), .ZN(prince_SR_Inv_Result_s2[32]) );
  XNOR2_X1 prince_AddKey2_XORInst_4_0_U1 ( .A(1'b0), .B(input_s2[16]), .ZN(
        prince_AddKey2_XORInst_4_0_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_4_1_U2 ( .A(prince_AddKey2_XORInst_4_1_n3), 
        .B(prince_selected_Key2_17_), .ZN(prince_SR_Inv_Result_s2[33]) );
  XNOR2_X1 prince_AddKey2_XORInst_4_1_U1 ( .A(1'b0), .B(input_s2[17]), .ZN(
        prince_AddKey2_XORInst_4_1_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_4_2_U2 ( .A(prince_AddKey2_XORInst_4_2_n3), 
        .B(prince_selected_Key2_18_), .ZN(prince_SR_Inv_Result_s2[34]) );
  XNOR2_X1 prince_AddKey2_XORInst_4_2_U1 ( .A(1'b0), .B(input_s2[18]), .ZN(
        prince_AddKey2_XORInst_4_2_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_4_3_U2 ( .A(prince_AddKey2_XORInst_4_3_n3), 
        .B(prince_selected_Key2_19_), .ZN(prince_SR_Inv_Result_s2[35]) );
  XNOR2_X1 prince_AddKey2_XORInst_4_3_U1 ( .A(1'b0), .B(input_s2[19]), .ZN(
        prince_AddKey2_XORInst_4_3_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_5_0_U2 ( .A(prince_AddKey2_XORInst_5_0_n3), 
        .B(prince_selected_Key2_20_), .ZN(prince_SR_Inv_Result_s2[52]) );
  XNOR2_X1 prince_AddKey2_XORInst_5_0_U1 ( .A(1'b0), .B(input_s2[20]), .ZN(
        prince_AddKey2_XORInst_5_0_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_5_1_U2 ( .A(prince_AddKey2_XORInst_5_1_n3), 
        .B(prince_selected_Key2_21_), .ZN(prince_SR_Inv_Result_s2[53]) );
  XNOR2_X1 prince_AddKey2_XORInst_5_1_U1 ( .A(1'b0), .B(input_s2[21]), .ZN(
        prince_AddKey2_XORInst_5_1_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_5_2_U2 ( .A(prince_AddKey2_XORInst_5_2_n3), 
        .B(prince_selected_Key2_22_), .ZN(prince_SR_Inv_Result_s2[54]) );
  XNOR2_X1 prince_AddKey2_XORInst_5_2_U1 ( .A(1'b0), .B(input_s2[22]), .ZN(
        prince_AddKey2_XORInst_5_2_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_5_3_U2 ( .A(prince_AddKey2_XORInst_5_3_n3), 
        .B(prince_selected_Key2_23_), .ZN(prince_SR_Inv_Result_s2[55]) );
  XNOR2_X1 prince_AddKey2_XORInst_5_3_U1 ( .A(1'b0), .B(input_s2[23]), .ZN(
        prince_AddKey2_XORInst_5_3_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_6_0_U2 ( .A(prince_AddKey2_XORInst_6_0_n3), 
        .B(prince_selected_Key2_24_), .ZN(prince_SR_Inv_Result_s2[8]) );
  XNOR2_X1 prince_AddKey2_XORInst_6_0_U1 ( .A(1'b0), .B(input_s2[24]), .ZN(
        prince_AddKey2_XORInst_6_0_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_6_1_U2 ( .A(prince_AddKey2_XORInst_6_1_n3), 
        .B(prince_selected_Key2_25_), .ZN(prince_SR_Inv_Result_s2[9]) );
  XNOR2_X1 prince_AddKey2_XORInst_6_1_U1 ( .A(1'b0), .B(input_s2[25]), .ZN(
        prince_AddKey2_XORInst_6_1_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_6_2_U2 ( .A(prince_AddKey2_XORInst_6_2_n3), 
        .B(prince_selected_Key2_26_), .ZN(prince_SR_Inv_Result_s2[10]) );
  XNOR2_X1 prince_AddKey2_XORInst_6_2_U1 ( .A(1'b0), .B(input_s2[26]), .ZN(
        prince_AddKey2_XORInst_6_2_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_6_3_U2 ( .A(prince_AddKey2_XORInst_6_3_n3), 
        .B(prince_selected_Key2_27_), .ZN(prince_SR_Inv_Result_s2[11]) );
  XNOR2_X1 prince_AddKey2_XORInst_6_3_U1 ( .A(1'b0), .B(input_s2[27]), .ZN(
        prince_AddKey2_XORInst_6_3_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_7_0_U2 ( .A(prince_AddKey2_XORInst_7_0_n3), 
        .B(prince_selected_Key2_28_), .ZN(prince_SR_Inv_Result_s2[28]) );
  XNOR2_X1 prince_AddKey2_XORInst_7_0_U1 ( .A(1'b0), .B(input_s2[28]), .ZN(
        prince_AddKey2_XORInst_7_0_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_7_1_U2 ( .A(prince_AddKey2_XORInst_7_1_n3), 
        .B(prince_selected_Key2_29_), .ZN(prince_SR_Inv_Result_s2[29]) );
  XNOR2_X1 prince_AddKey2_XORInst_7_1_U1 ( .A(1'b0), .B(input_s2[29]), .ZN(
        prince_AddKey2_XORInst_7_1_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_7_2_U2 ( .A(prince_AddKey2_XORInst_7_2_n3), 
        .B(prince_selected_Key2_30_), .ZN(prince_SR_Inv_Result_s2[30]) );
  XNOR2_X1 prince_AddKey2_XORInst_7_2_U1 ( .A(1'b0), .B(input_s2[30]), .ZN(
        prince_AddKey2_XORInst_7_2_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_7_3_U2 ( .A(prince_AddKey2_XORInst_7_3_n3), 
        .B(prince_selected_Key2_31_), .ZN(prince_SR_Inv_Result_s2[31]) );
  XNOR2_X1 prince_AddKey2_XORInst_7_3_U1 ( .A(1'b0), .B(input_s2[31]), .ZN(
        prince_AddKey2_XORInst_7_3_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_8_0_U2 ( .A(prince_AddKey2_XORInst_8_0_n3), 
        .B(prince_selected_Key2_32_), .ZN(prince_SR_Inv_Result_s2[48]) );
  XNOR2_X1 prince_AddKey2_XORInst_8_0_U1 ( .A(1'b0), .B(input_s2[32]), .ZN(
        prince_AddKey2_XORInst_8_0_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_8_1_U2 ( .A(prince_AddKey2_XORInst_8_1_n3), 
        .B(prince_selected_Key2_33_), .ZN(prince_SR_Inv_Result_s2[49]) );
  XNOR2_X1 prince_AddKey2_XORInst_8_1_U1 ( .A(1'b0), .B(input_s2[33]), .ZN(
        prince_AddKey2_XORInst_8_1_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_8_2_U2 ( .A(prince_AddKey2_XORInst_8_2_n3), 
        .B(prince_selected_Key2_34_), .ZN(prince_SR_Inv_Result_s2[50]) );
  XNOR2_X1 prince_AddKey2_XORInst_8_2_U1 ( .A(1'b0), .B(input_s2[34]), .ZN(
        prince_AddKey2_XORInst_8_2_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_8_3_U2 ( .A(prince_AddKey2_XORInst_8_3_n3), 
        .B(prince_selected_Key2_35_), .ZN(prince_SR_Inv_Result_s2[51]) );
  XNOR2_X1 prince_AddKey2_XORInst_8_3_U1 ( .A(1'b0), .B(input_s2[35]), .ZN(
        prince_AddKey2_XORInst_8_3_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_9_0_U2 ( .A(prince_AddKey2_XORInst_9_0_n3), 
        .B(prince_selected_Key2_36_), .ZN(prince_SR_Inv_Result_s2[4]) );
  XNOR2_X1 prince_AddKey2_XORInst_9_0_U1 ( .A(1'b0), .B(input_s2[36]), .ZN(
        prince_AddKey2_XORInst_9_0_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_9_1_U2 ( .A(prince_AddKey2_XORInst_9_1_n3), 
        .B(prince_selected_Key2_37_), .ZN(prince_SR_Inv_Result_s2[5]) );
  XNOR2_X1 prince_AddKey2_XORInst_9_1_U1 ( .A(1'b0), .B(input_s2[37]), .ZN(
        prince_AddKey2_XORInst_9_1_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_9_2_U2 ( .A(prince_AddKey2_XORInst_9_2_n3), 
        .B(prince_selected_Key2_38_), .ZN(prince_SR_Inv_Result_s2[6]) );
  XNOR2_X1 prince_AddKey2_XORInst_9_2_U1 ( .A(1'b0), .B(input_s2[38]), .ZN(
        prince_AddKey2_XORInst_9_2_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_9_3_U2 ( .A(prince_AddKey2_XORInst_9_3_n3), 
        .B(prince_selected_Key2_39_), .ZN(prince_SR_Inv_Result_s2[7]) );
  XNOR2_X1 prince_AddKey2_XORInst_9_3_U1 ( .A(1'b0), .B(input_s2[39]), .ZN(
        prince_AddKey2_XORInst_9_3_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_10_0_U2 ( .A(prince_AddKey2_XORInst_10_0_n3), 
        .B(prince_selected_Key2_40_), .ZN(prince_SR_Inv_Result_s2[24]) );
  XNOR2_X1 prince_AddKey2_XORInst_10_0_U1 ( .A(1'b0), .B(input_s2[40]), .ZN(
        prince_AddKey2_XORInst_10_0_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_10_1_U2 ( .A(prince_AddKey2_XORInst_10_1_n3), 
        .B(prince_selected_Key2_41_), .ZN(prince_SR_Inv_Result_s2[25]) );
  XNOR2_X1 prince_AddKey2_XORInst_10_1_U1 ( .A(1'b0), .B(input_s2[41]), .ZN(
        prince_AddKey2_XORInst_10_1_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_10_2_U2 ( .A(prince_AddKey2_XORInst_10_2_n3), 
        .B(prince_selected_Key2_42_), .ZN(prince_SR_Inv_Result_s2[26]) );
  XNOR2_X1 prince_AddKey2_XORInst_10_2_U1 ( .A(1'b0), .B(input_s2[42]), .ZN(
        prince_AddKey2_XORInst_10_2_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_10_3_U2 ( .A(prince_AddKey2_XORInst_10_3_n3), 
        .B(prince_selected_Key2_43_), .ZN(prince_SR_Inv_Result_s2[27]) );
  XNOR2_X1 prince_AddKey2_XORInst_10_3_U1 ( .A(1'b0), .B(input_s2[43]), .ZN(
        prince_AddKey2_XORInst_10_3_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_11_0_U2 ( .A(prince_AddKey2_XORInst_11_0_n3), 
        .B(prince_selected_Key2_44_), .ZN(prince_SR_Inv_Result_s2[44]) );
  XNOR2_X1 prince_AddKey2_XORInst_11_0_U1 ( .A(1'b0), .B(input_s2[44]), .ZN(
        prince_AddKey2_XORInst_11_0_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_11_1_U2 ( .A(prince_AddKey2_XORInst_11_1_n3), 
        .B(prince_selected_Key2_45_), .ZN(prince_SR_Inv_Result_s2[45]) );
  XNOR2_X1 prince_AddKey2_XORInst_11_1_U1 ( .A(1'b0), .B(input_s2[45]), .ZN(
        prince_AddKey2_XORInst_11_1_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_11_2_U2 ( .A(prince_AddKey2_XORInst_11_2_n3), 
        .B(prince_selected_Key2_46_), .ZN(prince_SR_Inv_Result_s2[46]) );
  XNOR2_X1 prince_AddKey2_XORInst_11_2_U1 ( .A(1'b0), .B(input_s2[46]), .ZN(
        prince_AddKey2_XORInst_11_2_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_11_3_U2 ( .A(prince_AddKey2_XORInst_11_3_n3), 
        .B(prince_selected_Key2_47_), .ZN(prince_SR_Inv_Result_s2[47]) );
  XNOR2_X1 prince_AddKey2_XORInst_11_3_U1 ( .A(1'b0), .B(input_s2[47]), .ZN(
        prince_AddKey2_XORInst_11_3_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_12_0_U2 ( .A(prince_AddKey2_XORInst_12_0_n3), 
        .B(prince_selected_Key2_48_), .ZN(prince_SR_Inv_Result_s2[0]) );
  XNOR2_X1 prince_AddKey2_XORInst_12_0_U1 ( .A(1'b0), .B(input_s2[48]), .ZN(
        prince_AddKey2_XORInst_12_0_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_12_1_U2 ( .A(prince_AddKey2_XORInst_12_1_n3), 
        .B(prince_selected_Key2_49_), .ZN(prince_SR_Inv_Result_s2[1]) );
  XNOR2_X1 prince_AddKey2_XORInst_12_1_U1 ( .A(1'b0), .B(input_s2[49]), .ZN(
        prince_AddKey2_XORInst_12_1_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_12_2_U2 ( .A(prince_AddKey2_XORInst_12_2_n3), 
        .B(prince_selected_Key2_50_), .ZN(prince_SR_Inv_Result_s2[2]) );
  XNOR2_X1 prince_AddKey2_XORInst_12_2_U1 ( .A(1'b0), .B(input_s2[50]), .ZN(
        prince_AddKey2_XORInst_12_2_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_12_3_U2 ( .A(prince_AddKey2_XORInst_12_3_n3), 
        .B(prince_selected_Key2_51_), .ZN(prince_SR_Inv_Result_s2[3]) );
  XNOR2_X1 prince_AddKey2_XORInst_12_3_U1 ( .A(1'b0), .B(input_s2[51]), .ZN(
        prince_AddKey2_XORInst_12_3_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_13_0_U2 ( .A(prince_AddKey2_XORInst_13_0_n3), 
        .B(prince_selected_Key2_52_), .ZN(prince_SR_Inv_Result_s2[20]) );
  XNOR2_X1 prince_AddKey2_XORInst_13_0_U1 ( .A(1'b0), .B(input_s2[52]), .ZN(
        prince_AddKey2_XORInst_13_0_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_13_1_U2 ( .A(prince_AddKey2_XORInst_13_1_n3), 
        .B(prince_selected_Key2_53_), .ZN(prince_SR_Inv_Result_s2[21]) );
  XNOR2_X1 prince_AddKey2_XORInst_13_1_U1 ( .A(1'b0), .B(input_s2[53]), .ZN(
        prince_AddKey2_XORInst_13_1_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_13_2_U2 ( .A(prince_AddKey2_XORInst_13_2_n3), 
        .B(prince_selected_Key2_54_), .ZN(prince_SR_Inv_Result_s2[22]) );
  XNOR2_X1 prince_AddKey2_XORInst_13_2_U1 ( .A(1'b0), .B(input_s2[54]), .ZN(
        prince_AddKey2_XORInst_13_2_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_13_3_U2 ( .A(prince_AddKey2_XORInst_13_3_n3), 
        .B(prince_selected_Key2_55_), .ZN(prince_SR_Inv_Result_s2[23]) );
  XNOR2_X1 prince_AddKey2_XORInst_13_3_U1 ( .A(1'b0), .B(input_s2[55]), .ZN(
        prince_AddKey2_XORInst_13_3_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_14_0_U2 ( .A(prince_AddKey2_XORInst_14_0_n3), 
        .B(prince_selected_Key2_56_), .ZN(prince_SR_Inv_Result_s2[40]) );
  XNOR2_X1 prince_AddKey2_XORInst_14_0_U1 ( .A(1'b0), .B(input_s2[56]), .ZN(
        prince_AddKey2_XORInst_14_0_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_14_1_U2 ( .A(prince_AddKey2_XORInst_14_1_n3), 
        .B(prince_selected_Key2_57_), .ZN(prince_SR_Inv_Result_s2[41]) );
  XNOR2_X1 prince_AddKey2_XORInst_14_1_U1 ( .A(1'b0), .B(input_s2[57]), .ZN(
        prince_AddKey2_XORInst_14_1_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_14_2_U2 ( .A(prince_AddKey2_XORInst_14_2_n3), 
        .B(prince_selected_Key2_58_), .ZN(prince_SR_Inv_Result_s2[42]) );
  XNOR2_X1 prince_AddKey2_XORInst_14_2_U1 ( .A(1'b0), .B(input_s2[58]), .ZN(
        prince_AddKey2_XORInst_14_2_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_14_3_U2 ( .A(prince_AddKey2_XORInst_14_3_n3), 
        .B(prince_selected_Key2_59_), .ZN(prince_SR_Inv_Result_s2[43]) );
  XNOR2_X1 prince_AddKey2_XORInst_14_3_U1 ( .A(1'b0), .B(input_s2[59]), .ZN(
        prince_AddKey2_XORInst_14_3_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_15_0_U2 ( .A(prince_AddKey2_XORInst_15_0_n3), 
        .B(prince_selected_Key2_60_), .ZN(prince_SR_Inv_Result_s2[60]) );
  XNOR2_X1 prince_AddKey2_XORInst_15_0_U1 ( .A(1'b0), .B(input_s2[60]), .ZN(
        prince_AddKey2_XORInst_15_0_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_15_1_U2 ( .A(prince_AddKey2_XORInst_15_1_n3), 
        .B(prince_selected_Key2_61_), .ZN(prince_SR_Inv_Result_s2[61]) );
  XNOR2_X1 prince_AddKey2_XORInst_15_1_U1 ( .A(1'b0), .B(input_s2[61]), .ZN(
        prince_AddKey2_XORInst_15_1_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_15_2_U2 ( .A(prince_AddKey2_XORInst_15_2_n3), 
        .B(prince_selected_Key2_62_), .ZN(prince_SR_Inv_Result_s2[62]) );
  XNOR2_X1 prince_AddKey2_XORInst_15_2_U1 ( .A(1'b0), .B(input_s2[62]), .ZN(
        prince_AddKey2_XORInst_15_2_n3) );
  XNOR2_X1 prince_AddKey2_XORInst_15_3_U2 ( .A(prince_AddKey2_XORInst_15_3_n3), 
        .B(prince_selected_Key2_63_), .ZN(prince_SR_Inv_Result_s2[63]) );
  XNOR2_X1 prince_AddKey2_XORInst_15_3_U1 ( .A(1'b0), .B(input_s2[63]), .ZN(
        prince_AddKey2_XORInst_15_3_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_0_0_U2 ( .A(prince_AddKey3_XORInst_0_0_n3), 
        .B(prince_selected_Key3_0_), .ZN(prince_SR_Inv_Result_s3[16]) );
  XNOR2_X1 prince_AddKey3_XORInst_0_0_U1 ( .A(1'b0), .B(input_s3[0]), .ZN(
        prince_AddKey3_XORInst_0_0_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_0_1_U2 ( .A(prince_AddKey3_XORInst_0_1_n3), 
        .B(prince_selected_Key3_1_), .ZN(prince_SR_Inv_Result_s3[17]) );
  XNOR2_X1 prince_AddKey3_XORInst_0_1_U1 ( .A(1'b0), .B(input_s3[1]), .ZN(
        prince_AddKey3_XORInst_0_1_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_0_2_U2 ( .A(prince_AddKey3_XORInst_0_2_n3), 
        .B(prince_selected_Key3_2_), .ZN(prince_SR_Inv_Result_s3[18]) );
  XNOR2_X1 prince_AddKey3_XORInst_0_2_U1 ( .A(1'b0), .B(input_s3[2]), .ZN(
        prince_AddKey3_XORInst_0_2_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_0_3_U2 ( .A(prince_AddKey3_XORInst_0_3_n3), 
        .B(prince_selected_Key3_3_), .ZN(prince_SR_Inv_Result_s3[19]) );
  XNOR2_X1 prince_AddKey3_XORInst_0_3_U1 ( .A(1'b0), .B(input_s3[3]), .ZN(
        prince_AddKey3_XORInst_0_3_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_1_0_U2 ( .A(prince_AddKey3_XORInst_1_0_n3), 
        .B(prince_selected_Key3_4_), .ZN(prince_SR_Inv_Result_s3[36]) );
  XNOR2_X1 prince_AddKey3_XORInst_1_0_U1 ( .A(1'b0), .B(input_s3[4]), .ZN(
        prince_AddKey3_XORInst_1_0_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_1_1_U2 ( .A(prince_AddKey3_XORInst_1_1_n3), 
        .B(prince_selected_Key3_5_), .ZN(prince_SR_Inv_Result_s3[37]) );
  XNOR2_X1 prince_AddKey3_XORInst_1_1_U1 ( .A(1'b0), .B(input_s3[5]), .ZN(
        prince_AddKey3_XORInst_1_1_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_1_2_U2 ( .A(prince_AddKey3_XORInst_1_2_n3), 
        .B(prince_selected_Key3_6_), .ZN(prince_SR_Inv_Result_s3[38]) );
  XNOR2_X1 prince_AddKey3_XORInst_1_2_U1 ( .A(1'b0), .B(input_s3[6]), .ZN(
        prince_AddKey3_XORInst_1_2_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_1_3_U2 ( .A(prince_AddKey3_XORInst_1_3_n3), 
        .B(prince_selected_Key3_7_), .ZN(prince_SR_Inv_Result_s3[39]) );
  XNOR2_X1 prince_AddKey3_XORInst_1_3_U1 ( .A(1'b0), .B(input_s3[7]), .ZN(
        prince_AddKey3_XORInst_1_3_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_2_0_U2 ( .A(prince_AddKey3_XORInst_2_0_n3), 
        .B(prince_selected_Key3_8_), .ZN(prince_SR_Inv_Result_s3[56]) );
  XNOR2_X1 prince_AddKey3_XORInst_2_0_U1 ( .A(1'b0), .B(input_s3[8]), .ZN(
        prince_AddKey3_XORInst_2_0_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_2_1_U2 ( .A(prince_AddKey3_XORInst_2_1_n3), 
        .B(prince_selected_Key3_9_), .ZN(prince_SR_Inv_Result_s3[57]) );
  XNOR2_X1 prince_AddKey3_XORInst_2_1_U1 ( .A(1'b0), .B(input_s3[9]), .ZN(
        prince_AddKey3_XORInst_2_1_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_2_2_U2 ( .A(prince_AddKey3_XORInst_2_2_n3), 
        .B(prince_selected_Key3_10_), .ZN(prince_SR_Inv_Result_s3[58]) );
  XNOR2_X1 prince_AddKey3_XORInst_2_2_U1 ( .A(1'b0), .B(input_s3[10]), .ZN(
        prince_AddKey3_XORInst_2_2_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_2_3_U2 ( .A(prince_AddKey3_XORInst_2_3_n3), 
        .B(prince_selected_Key3_11_), .ZN(prince_SR_Inv_Result_s3[59]) );
  XNOR2_X1 prince_AddKey3_XORInst_2_3_U1 ( .A(1'b0), .B(input_s3[11]), .ZN(
        prince_AddKey3_XORInst_2_3_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_3_0_U2 ( .A(prince_AddKey3_XORInst_3_0_n3), 
        .B(prince_selected_Key3_12_), .ZN(prince_SR_Inv_Result_s3[12]) );
  XNOR2_X1 prince_AddKey3_XORInst_3_0_U1 ( .A(1'b0), .B(input_s3[12]), .ZN(
        prince_AddKey3_XORInst_3_0_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_3_1_U2 ( .A(prince_AddKey3_XORInst_3_1_n3), 
        .B(prince_selected_Key3_13_), .ZN(prince_SR_Inv_Result_s3[13]) );
  XNOR2_X1 prince_AddKey3_XORInst_3_1_U1 ( .A(1'b0), .B(input_s3[13]), .ZN(
        prince_AddKey3_XORInst_3_1_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_3_2_U2 ( .A(prince_AddKey3_XORInst_3_2_n3), 
        .B(prince_selected_Key3_14_), .ZN(prince_SR_Inv_Result_s3[14]) );
  XNOR2_X1 prince_AddKey3_XORInst_3_2_U1 ( .A(1'b0), .B(input_s3[14]), .ZN(
        prince_AddKey3_XORInst_3_2_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_3_3_U2 ( .A(prince_AddKey3_XORInst_3_3_n3), 
        .B(prince_selected_Key3_15_), .ZN(prince_SR_Inv_Result_s3[15]) );
  XNOR2_X1 prince_AddKey3_XORInst_3_3_U1 ( .A(1'b0), .B(input_s3[15]), .ZN(
        prince_AddKey3_XORInst_3_3_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_4_0_U2 ( .A(prince_AddKey3_XORInst_4_0_n3), 
        .B(prince_selected_Key3_16_), .ZN(prince_SR_Inv_Result_s3[32]) );
  XNOR2_X1 prince_AddKey3_XORInst_4_0_U1 ( .A(1'b0), .B(input_s3[16]), .ZN(
        prince_AddKey3_XORInst_4_0_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_4_1_U2 ( .A(prince_AddKey3_XORInst_4_1_n3), 
        .B(prince_selected_Key3_17_), .ZN(prince_SR_Inv_Result_s3[33]) );
  XNOR2_X1 prince_AddKey3_XORInst_4_1_U1 ( .A(1'b0), .B(input_s3[17]), .ZN(
        prince_AddKey3_XORInst_4_1_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_4_2_U2 ( .A(prince_AddKey3_XORInst_4_2_n3), 
        .B(prince_selected_Key3_18_), .ZN(prince_SR_Inv_Result_s3[34]) );
  XNOR2_X1 prince_AddKey3_XORInst_4_2_U1 ( .A(1'b0), .B(input_s3[18]), .ZN(
        prince_AddKey3_XORInst_4_2_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_4_3_U2 ( .A(prince_AddKey3_XORInst_4_3_n3), 
        .B(prince_selected_Key3_19_), .ZN(prince_SR_Inv_Result_s3[35]) );
  XNOR2_X1 prince_AddKey3_XORInst_4_3_U1 ( .A(1'b0), .B(input_s3[19]), .ZN(
        prince_AddKey3_XORInst_4_3_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_5_0_U2 ( .A(prince_AddKey3_XORInst_5_0_n3), 
        .B(prince_selected_Key3_20_), .ZN(prince_SR_Inv_Result_s3[52]) );
  XNOR2_X1 prince_AddKey3_XORInst_5_0_U1 ( .A(1'b0), .B(input_s3[20]), .ZN(
        prince_AddKey3_XORInst_5_0_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_5_1_U2 ( .A(prince_AddKey3_XORInst_5_1_n3), 
        .B(prince_selected_Key3_21_), .ZN(prince_SR_Inv_Result_s3[53]) );
  XNOR2_X1 prince_AddKey3_XORInst_5_1_U1 ( .A(1'b0), .B(input_s3[21]), .ZN(
        prince_AddKey3_XORInst_5_1_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_5_2_U2 ( .A(prince_AddKey3_XORInst_5_2_n3), 
        .B(prince_selected_Key3_22_), .ZN(prince_SR_Inv_Result_s3[54]) );
  XNOR2_X1 prince_AddKey3_XORInst_5_2_U1 ( .A(1'b0), .B(input_s3[22]), .ZN(
        prince_AddKey3_XORInst_5_2_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_5_3_U2 ( .A(prince_AddKey3_XORInst_5_3_n3), 
        .B(prince_selected_Key3_23_), .ZN(prince_SR_Inv_Result_s3[55]) );
  XNOR2_X1 prince_AddKey3_XORInst_5_3_U1 ( .A(1'b0), .B(input_s3[23]), .ZN(
        prince_AddKey3_XORInst_5_3_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_6_0_U2 ( .A(prince_AddKey3_XORInst_6_0_n3), 
        .B(prince_selected_Key3_24_), .ZN(prince_SR_Inv_Result_s3[8]) );
  XNOR2_X1 prince_AddKey3_XORInst_6_0_U1 ( .A(1'b0), .B(input_s3[24]), .ZN(
        prince_AddKey3_XORInst_6_0_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_6_1_U2 ( .A(prince_AddKey3_XORInst_6_1_n3), 
        .B(prince_selected_Key3_25_), .ZN(prince_SR_Inv_Result_s3[9]) );
  XNOR2_X1 prince_AddKey3_XORInst_6_1_U1 ( .A(1'b0), .B(input_s3[25]), .ZN(
        prince_AddKey3_XORInst_6_1_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_6_2_U2 ( .A(prince_AddKey3_XORInst_6_2_n3), 
        .B(prince_selected_Key3_26_), .ZN(prince_SR_Inv_Result_s3[10]) );
  XNOR2_X1 prince_AddKey3_XORInst_6_2_U1 ( .A(1'b0), .B(input_s3[26]), .ZN(
        prince_AddKey3_XORInst_6_2_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_6_3_U2 ( .A(prince_AddKey3_XORInst_6_3_n3), 
        .B(prince_selected_Key3_27_), .ZN(prince_SR_Inv_Result_s3[11]) );
  XNOR2_X1 prince_AddKey3_XORInst_6_3_U1 ( .A(1'b0), .B(input_s3[27]), .ZN(
        prince_AddKey3_XORInst_6_3_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_7_0_U2 ( .A(prince_AddKey3_XORInst_7_0_n3), 
        .B(prince_selected_Key3_28_), .ZN(prince_SR_Inv_Result_s3[28]) );
  XNOR2_X1 prince_AddKey3_XORInst_7_0_U1 ( .A(1'b0), .B(input_s3[28]), .ZN(
        prince_AddKey3_XORInst_7_0_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_7_1_U2 ( .A(prince_AddKey3_XORInst_7_1_n3), 
        .B(prince_selected_Key3_29_), .ZN(prince_SR_Inv_Result_s3[29]) );
  XNOR2_X1 prince_AddKey3_XORInst_7_1_U1 ( .A(1'b0), .B(input_s3[29]), .ZN(
        prince_AddKey3_XORInst_7_1_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_7_2_U2 ( .A(prince_AddKey3_XORInst_7_2_n3), 
        .B(prince_selected_Key3_30_), .ZN(prince_SR_Inv_Result_s3[30]) );
  XNOR2_X1 prince_AddKey3_XORInst_7_2_U1 ( .A(1'b0), .B(input_s3[30]), .ZN(
        prince_AddKey3_XORInst_7_2_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_7_3_U2 ( .A(prince_AddKey3_XORInst_7_3_n3), 
        .B(prince_selected_Key3_31_), .ZN(prince_SR_Inv_Result_s3[31]) );
  XNOR2_X1 prince_AddKey3_XORInst_7_3_U1 ( .A(1'b0), .B(input_s3[31]), .ZN(
        prince_AddKey3_XORInst_7_3_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_8_0_U2 ( .A(prince_AddKey3_XORInst_8_0_n3), 
        .B(prince_selected_Key3_32_), .ZN(prince_SR_Inv_Result_s3[48]) );
  XNOR2_X1 prince_AddKey3_XORInst_8_0_U1 ( .A(1'b0), .B(input_s3[32]), .ZN(
        prince_AddKey3_XORInst_8_0_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_8_1_U2 ( .A(prince_AddKey3_XORInst_8_1_n3), 
        .B(prince_selected_Key3_33_), .ZN(prince_SR_Inv_Result_s3[49]) );
  XNOR2_X1 prince_AddKey3_XORInst_8_1_U1 ( .A(1'b0), .B(input_s3[33]), .ZN(
        prince_AddKey3_XORInst_8_1_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_8_2_U2 ( .A(prince_AddKey3_XORInst_8_2_n3), 
        .B(prince_selected_Key3_34_), .ZN(prince_SR_Inv_Result_s3[50]) );
  XNOR2_X1 prince_AddKey3_XORInst_8_2_U1 ( .A(1'b0), .B(input_s3[34]), .ZN(
        prince_AddKey3_XORInst_8_2_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_8_3_U2 ( .A(prince_AddKey3_XORInst_8_3_n3), 
        .B(prince_selected_Key3_35_), .ZN(prince_SR_Inv_Result_s3[51]) );
  XNOR2_X1 prince_AddKey3_XORInst_8_3_U1 ( .A(1'b0), .B(input_s3[35]), .ZN(
        prince_AddKey3_XORInst_8_3_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_9_0_U2 ( .A(prince_AddKey3_XORInst_9_0_n3), 
        .B(prince_selected_Key3_36_), .ZN(prince_SR_Inv_Result_s3[4]) );
  XNOR2_X1 prince_AddKey3_XORInst_9_0_U1 ( .A(1'b0), .B(input_s3[36]), .ZN(
        prince_AddKey3_XORInst_9_0_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_9_1_U2 ( .A(prince_AddKey3_XORInst_9_1_n3), 
        .B(prince_selected_Key3_37_), .ZN(prince_SR_Inv_Result_s3[5]) );
  XNOR2_X1 prince_AddKey3_XORInst_9_1_U1 ( .A(1'b0), .B(input_s3[37]), .ZN(
        prince_AddKey3_XORInst_9_1_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_9_2_U2 ( .A(prince_AddKey3_XORInst_9_2_n3), 
        .B(prince_selected_Key3_38_), .ZN(prince_SR_Inv_Result_s3[6]) );
  XNOR2_X1 prince_AddKey3_XORInst_9_2_U1 ( .A(1'b0), .B(input_s3[38]), .ZN(
        prince_AddKey3_XORInst_9_2_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_9_3_U2 ( .A(prince_AddKey3_XORInst_9_3_n3), 
        .B(prince_selected_Key3_39_), .ZN(prince_SR_Inv_Result_s3[7]) );
  XNOR2_X1 prince_AddKey3_XORInst_9_3_U1 ( .A(1'b0), .B(input_s3[39]), .ZN(
        prince_AddKey3_XORInst_9_3_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_10_0_U2 ( .A(prince_AddKey3_XORInst_10_0_n3), 
        .B(prince_selected_Key3_40_), .ZN(prince_SR_Inv_Result_s3[24]) );
  XNOR2_X1 prince_AddKey3_XORInst_10_0_U1 ( .A(1'b0), .B(input_s3[40]), .ZN(
        prince_AddKey3_XORInst_10_0_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_10_1_U2 ( .A(prince_AddKey3_XORInst_10_1_n3), 
        .B(prince_selected_Key3_41_), .ZN(prince_SR_Inv_Result_s3[25]) );
  XNOR2_X1 prince_AddKey3_XORInst_10_1_U1 ( .A(1'b0), .B(input_s3[41]), .ZN(
        prince_AddKey3_XORInst_10_1_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_10_2_U2 ( .A(prince_AddKey3_XORInst_10_2_n3), 
        .B(prince_selected_Key3_42_), .ZN(prince_SR_Inv_Result_s3[26]) );
  XNOR2_X1 prince_AddKey3_XORInst_10_2_U1 ( .A(1'b0), .B(input_s3[42]), .ZN(
        prince_AddKey3_XORInst_10_2_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_10_3_U2 ( .A(prince_AddKey3_XORInst_10_3_n3), 
        .B(prince_selected_Key3_43_), .ZN(prince_SR_Inv_Result_s3[27]) );
  XNOR2_X1 prince_AddKey3_XORInst_10_3_U1 ( .A(1'b0), .B(input_s3[43]), .ZN(
        prince_AddKey3_XORInst_10_3_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_11_0_U2 ( .A(prince_AddKey3_XORInst_11_0_n3), 
        .B(prince_selected_Key3_44_), .ZN(prince_SR_Inv_Result_s3[44]) );
  XNOR2_X1 prince_AddKey3_XORInst_11_0_U1 ( .A(1'b0), .B(input_s3[44]), .ZN(
        prince_AddKey3_XORInst_11_0_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_11_1_U2 ( .A(prince_AddKey3_XORInst_11_1_n3), 
        .B(prince_selected_Key3_45_), .ZN(prince_SR_Inv_Result_s3[45]) );
  XNOR2_X1 prince_AddKey3_XORInst_11_1_U1 ( .A(1'b0), .B(input_s3[45]), .ZN(
        prince_AddKey3_XORInst_11_1_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_11_2_U2 ( .A(prince_AddKey3_XORInst_11_2_n3), 
        .B(prince_selected_Key3_46_), .ZN(prince_SR_Inv_Result_s3[46]) );
  XNOR2_X1 prince_AddKey3_XORInst_11_2_U1 ( .A(1'b0), .B(input_s3[46]), .ZN(
        prince_AddKey3_XORInst_11_2_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_11_3_U2 ( .A(prince_AddKey3_XORInst_11_3_n3), 
        .B(prince_selected_Key3_47_), .ZN(prince_SR_Inv_Result_s3[47]) );
  XNOR2_X1 prince_AddKey3_XORInst_11_3_U1 ( .A(1'b0), .B(input_s3[47]), .ZN(
        prince_AddKey3_XORInst_11_3_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_12_0_U2 ( .A(prince_AddKey3_XORInst_12_0_n3), 
        .B(prince_selected_Key3_48_), .ZN(prince_SR_Inv_Result_s3[0]) );
  XNOR2_X1 prince_AddKey3_XORInst_12_0_U1 ( .A(1'b0), .B(input_s3[48]), .ZN(
        prince_AddKey3_XORInst_12_0_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_12_1_U2 ( .A(prince_AddKey3_XORInst_12_1_n3), 
        .B(prince_selected_Key3_49_), .ZN(prince_SR_Inv_Result_s3[1]) );
  XNOR2_X1 prince_AddKey3_XORInst_12_1_U1 ( .A(1'b0), .B(input_s3[49]), .ZN(
        prince_AddKey3_XORInst_12_1_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_12_2_U2 ( .A(prince_AddKey3_XORInst_12_2_n3), 
        .B(prince_selected_Key3_50_), .ZN(prince_SR_Inv_Result_s3[2]) );
  XNOR2_X1 prince_AddKey3_XORInst_12_2_U1 ( .A(1'b0), .B(input_s3[50]), .ZN(
        prince_AddKey3_XORInst_12_2_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_12_3_U2 ( .A(prince_AddKey3_XORInst_12_3_n3), 
        .B(prince_selected_Key3_51_), .ZN(prince_SR_Inv_Result_s3[3]) );
  XNOR2_X1 prince_AddKey3_XORInst_12_3_U1 ( .A(1'b0), .B(input_s3[51]), .ZN(
        prince_AddKey3_XORInst_12_3_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_13_0_U2 ( .A(prince_AddKey3_XORInst_13_0_n3), 
        .B(prince_selected_Key3_52_), .ZN(prince_SR_Inv_Result_s3[20]) );
  XNOR2_X1 prince_AddKey3_XORInst_13_0_U1 ( .A(1'b0), .B(input_s3[52]), .ZN(
        prince_AddKey3_XORInst_13_0_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_13_1_U2 ( .A(prince_AddKey3_XORInst_13_1_n3), 
        .B(prince_selected_Key3_53_), .ZN(prince_SR_Inv_Result_s3[21]) );
  XNOR2_X1 prince_AddKey3_XORInst_13_1_U1 ( .A(1'b0), .B(input_s3[53]), .ZN(
        prince_AddKey3_XORInst_13_1_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_13_2_U2 ( .A(prince_AddKey3_XORInst_13_2_n3), 
        .B(prince_selected_Key3_54_), .ZN(prince_SR_Inv_Result_s3[22]) );
  XNOR2_X1 prince_AddKey3_XORInst_13_2_U1 ( .A(1'b0), .B(input_s3[54]), .ZN(
        prince_AddKey3_XORInst_13_2_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_13_3_U2 ( .A(prince_AddKey3_XORInst_13_3_n3), 
        .B(prince_selected_Key3_55_), .ZN(prince_SR_Inv_Result_s3[23]) );
  XNOR2_X1 prince_AddKey3_XORInst_13_3_U1 ( .A(1'b0), .B(input_s3[55]), .ZN(
        prince_AddKey3_XORInst_13_3_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_14_0_U2 ( .A(prince_AddKey3_XORInst_14_0_n3), 
        .B(prince_selected_Key3_56_), .ZN(prince_SR_Inv_Result_s3[40]) );
  XNOR2_X1 prince_AddKey3_XORInst_14_0_U1 ( .A(1'b0), .B(input_s3[56]), .ZN(
        prince_AddKey3_XORInst_14_0_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_14_1_U2 ( .A(prince_AddKey3_XORInst_14_1_n3), 
        .B(prince_selected_Key3_57_), .ZN(prince_SR_Inv_Result_s3[41]) );
  XNOR2_X1 prince_AddKey3_XORInst_14_1_U1 ( .A(1'b0), .B(input_s3[57]), .ZN(
        prince_AddKey3_XORInst_14_1_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_14_2_U2 ( .A(prince_AddKey3_XORInst_14_2_n3), 
        .B(prince_selected_Key3_58_), .ZN(prince_SR_Inv_Result_s3[42]) );
  XNOR2_X1 prince_AddKey3_XORInst_14_2_U1 ( .A(1'b0), .B(input_s3[58]), .ZN(
        prince_AddKey3_XORInst_14_2_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_14_3_U2 ( .A(prince_AddKey3_XORInst_14_3_n3), 
        .B(prince_selected_Key3_59_), .ZN(prince_SR_Inv_Result_s3[43]) );
  XNOR2_X1 prince_AddKey3_XORInst_14_3_U1 ( .A(1'b0), .B(input_s3[59]), .ZN(
        prince_AddKey3_XORInst_14_3_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_15_0_U2 ( .A(prince_AddKey3_XORInst_15_0_n3), 
        .B(prince_selected_Key3_60_), .ZN(prince_SR_Inv_Result_s3[60]) );
  XNOR2_X1 prince_AddKey3_XORInst_15_0_U1 ( .A(1'b0), .B(input_s3[60]), .ZN(
        prince_AddKey3_XORInst_15_0_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_15_1_U2 ( .A(prince_AddKey3_XORInst_15_1_n3), 
        .B(prince_selected_Key3_61_), .ZN(prince_SR_Inv_Result_s3[61]) );
  XNOR2_X1 prince_AddKey3_XORInst_15_1_U1 ( .A(1'b0), .B(input_s3[61]), .ZN(
        prince_AddKey3_XORInst_15_1_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_15_2_U2 ( .A(prince_AddKey3_XORInst_15_2_n3), 
        .B(prince_selected_Key3_62_), .ZN(prince_SR_Inv_Result_s3[62]) );
  XNOR2_X1 prince_AddKey3_XORInst_15_2_U1 ( .A(1'b0), .B(input_s3[62]), .ZN(
        prince_AddKey3_XORInst_15_2_n3) );
  XNOR2_X1 prince_AddKey3_XORInst_15_3_U2 ( .A(prince_AddKey3_XORInst_15_3_n3), 
        .B(prince_selected_Key3_63_), .ZN(prince_SR_Inv_Result_s3[63]) );
  XNOR2_X1 prince_AddKey3_XORInst_15_3_U1 ( .A(1'b0), .B(input_s3[63]), .ZN(
        prince_AddKey3_XORInst_15_3_n3) );
  XNOR2_X1 prince_rounds_U241 ( .A(prince_rounds_SR_Inv_Result_s3[57]), .B(
        prince_rounds_n65), .ZN(prince_rounds_Output_s3[9]) );
  XNOR2_X1 prince_rounds_U240 ( .A(prince_rounds_SR_Inv_Result_s3[56]), .B(
        prince_rounds_n64), .ZN(prince_rounds_Output_s3[8]) );
  XNOR2_X1 prince_rounds_U239 ( .A(prince_rounds_SR_Inv_Result_s3[39]), .B(
        prince_rounds_n63), .ZN(prince_rounds_Output_s3[7]) );
  XNOR2_X1 prince_rounds_U238 ( .A(prince_rounds_SR_Inv_Result_s3[38]), .B(
        prince_rounds_n62), .ZN(prince_rounds_Output_s3[6]) );
  XNOR2_X1 prince_rounds_U237 ( .A(prince_rounds_SR_Inv_Result_s3[63]), .B(
        prince_rounds_n61), .ZN(prince_rounds_Output_s3[63]) );
  XNOR2_X1 prince_rounds_U236 ( .A(prince_rounds_SR_Inv_Result_s3[62]), .B(
        prince_rounds_n60), .ZN(prince_rounds_Output_s3[62]) );
  XNOR2_X1 prince_rounds_U235 ( .A(prince_rounds_SR_Inv_Result_s3[61]), .B(
        prince_rounds_n59), .ZN(prince_rounds_Output_s3[61]) );
  XNOR2_X1 prince_rounds_U234 ( .A(prince_rounds_SR_Inv_Result_s3[60]), .B(
        prince_rounds_n58), .ZN(prince_rounds_Output_s3[60]) );
  XNOR2_X1 prince_rounds_U233 ( .A(prince_rounds_SR_Inv_Result_s3[37]), .B(
        prince_rounds_n57), .ZN(prince_rounds_Output_s3[5]) );
  XNOR2_X1 prince_rounds_U232 ( .A(prince_rounds_SR_Inv_Result_s3[43]), .B(
        prince_rounds_n56), .ZN(prince_rounds_Output_s3[59]) );
  XNOR2_X1 prince_rounds_U231 ( .A(prince_rounds_SR_Inv_Result_s3[42]), .B(
        prince_rounds_n55), .ZN(prince_rounds_Output_s3[58]) );
  XNOR2_X1 prince_rounds_U230 ( .A(prince_rounds_SR_Inv_Result_s3[41]), .B(
        prince_rounds_n65), .ZN(prince_rounds_Output_s3[57]) );
  XNOR2_X1 prince_rounds_U229 ( .A(prince_rounds_SR_Inv_Result_s3[40]), .B(
        prince_rounds_n64), .ZN(prince_rounds_Output_s3[56]) );
  XNOR2_X1 prince_rounds_U228 ( .A(prince_rounds_SR_Inv_Result_s3[23]), .B(
        prince_rounds_n63), .ZN(prince_rounds_Output_s3[55]) );
  XNOR2_X1 prince_rounds_U227 ( .A(prince_rounds_SR_Inv_Result_s3[22]), .B(
        prince_rounds_n62), .ZN(prince_rounds_Output_s3[54]) );
  XNOR2_X1 prince_rounds_U226 ( .A(prince_rounds_SR_Inv_Result_s3[21]), .B(
        prince_rounds_n57), .ZN(prince_rounds_Output_s3[53]) );
  XNOR2_X1 prince_rounds_U225 ( .A(prince_rounds_SR_Inv_Result_s3[20]), .B(
        prince_rounds_n54), .ZN(prince_rounds_Output_s3[52]) );
  XNOR2_X1 prince_rounds_U224 ( .A(prince_rounds_SR_Inv_Result_s3[3]), .B(
        prince_rounds_n53), .ZN(prince_rounds_Output_s3[51]) );
  XNOR2_X1 prince_rounds_U223 ( .A(prince_rounds_SR_Inv_Result_s3[2]), .B(
        prince_rounds_n52), .ZN(prince_rounds_Output_s3[50]) );
  XNOR2_X1 prince_rounds_U222 ( .A(prince_rounds_SR_Inv_Result_s3[36]), .B(
        prince_rounds_n54), .ZN(prince_rounds_Output_s3[4]) );
  XNOR2_X1 prince_rounds_U221 ( .A(prince_rounds_SR_Inv_Result_s3[1]), .B(
        prince_rounds_n51), .ZN(prince_rounds_Output_s3[49]) );
  XNOR2_X1 prince_rounds_U220 ( .A(prince_rounds_SR_Inv_Result_s3[0]), .B(
        prince_rounds_n50), .ZN(prince_rounds_Output_s3[48]) );
  XNOR2_X1 prince_rounds_U219 ( .A(prince_rounds_SR_Inv_Result_s3[47]), .B(
        prince_rounds_n61), .ZN(prince_rounds_Output_s3[47]) );
  XNOR2_X1 prince_rounds_U218 ( .A(prince_rounds_SR_Inv_Result_s3[46]), .B(
        prince_rounds_n60), .ZN(prince_rounds_Output_s3[46]) );
  XNOR2_X1 prince_rounds_U217 ( .A(prince_rounds_SR_Inv_Result_s3[45]), .B(
        prince_rounds_n59), .ZN(prince_rounds_Output_s3[45]) );
  XNOR2_X1 prince_rounds_U216 ( .A(prince_rounds_SR_Inv_Result_s3[44]), .B(
        prince_rounds_n58), .ZN(prince_rounds_Output_s3[44]) );
  XNOR2_X1 prince_rounds_U215 ( .A(prince_rounds_SR_Inv_Result_s3[27]), .B(
        prince_rounds_n56), .ZN(prince_rounds_Output_s3[43]) );
  XNOR2_X1 prince_rounds_U214 ( .A(prince_rounds_SR_Inv_Result_s3[26]), .B(
        prince_rounds_n55), .ZN(prince_rounds_Output_s3[42]) );
  XNOR2_X1 prince_rounds_U213 ( .A(prince_rounds_SR_Inv_Result_s3[25]), .B(
        prince_rounds_n65), .ZN(prince_rounds_Output_s3[41]) );
  XNOR2_X1 prince_rounds_U212 ( .A(prince_rounds_SR_Inv_Result_s3[24]), .B(
        prince_rounds_n64), .ZN(prince_rounds_Output_s3[40]) );
  XNOR2_X1 prince_rounds_U211 ( .A(prince_rounds_SR_Inv_Result_s3[19]), .B(
        prince_rounds_n53), .ZN(prince_rounds_Output_s3[3]) );
  XNOR2_X1 prince_rounds_U210 ( .A(prince_rounds_SR_Inv_Result_s3[7]), .B(
        prince_rounds_n63), .ZN(prince_rounds_Output_s3[39]) );
  XNOR2_X1 prince_rounds_U209 ( .A(prince_rounds_SR_Inv_Result_s3[6]), .B(
        prince_rounds_n62), .ZN(prince_rounds_Output_s3[38]) );
  XNOR2_X1 prince_rounds_U208 ( .A(prince_rounds_SR_Inv_Result_s3[5]), .B(
        prince_rounds_n57), .ZN(prince_rounds_Output_s3[37]) );
  XNOR2_X1 prince_rounds_U207 ( .A(prince_rounds_SR_Inv_Result_s3[4]), .B(
        prince_rounds_n54), .ZN(prince_rounds_Output_s3[36]) );
  XNOR2_X1 prince_rounds_U206 ( .A(prince_rounds_SR_Inv_Result_s3[51]), .B(
        prince_rounds_n53), .ZN(prince_rounds_Output_s3[35]) );
  XNOR2_X1 prince_rounds_U205 ( .A(prince_rounds_SR_Inv_Result_s3[50]), .B(
        prince_rounds_n52), .ZN(prince_rounds_Output_s3[34]) );
  XNOR2_X1 prince_rounds_U204 ( .A(prince_rounds_SR_Inv_Result_s3[49]), .B(
        prince_rounds_n51), .ZN(prince_rounds_Output_s3[33]) );
  XNOR2_X1 prince_rounds_U203 ( .A(prince_rounds_SR_Inv_Result_s3[48]), .B(
        prince_rounds_n50), .ZN(prince_rounds_Output_s3[32]) );
  XNOR2_X1 prince_rounds_U202 ( .A(prince_rounds_SR_Inv_Result_s3[31]), .B(
        prince_rounds_n61), .ZN(prince_rounds_Output_s3[31]) );
  XNOR2_X1 prince_rounds_U201 ( .A(prince_rounds_SR_Inv_Result_s3[30]), .B(
        prince_rounds_n60), .ZN(prince_rounds_Output_s3[30]) );
  XNOR2_X1 prince_rounds_U200 ( .A(prince_rounds_SR_Inv_Result_s3[18]), .B(
        prince_rounds_n52), .ZN(prince_rounds_Output_s3[2]) );
  XNOR2_X1 prince_rounds_U199 ( .A(prince_rounds_SR_Inv_Result_s3[29]), .B(
        prince_rounds_n59), .ZN(prince_rounds_Output_s3[29]) );
  XNOR2_X1 prince_rounds_U198 ( .A(prince_rounds_SR_Inv_Result_s3[28]), .B(
        prince_rounds_n58), .ZN(prince_rounds_Output_s3[28]) );
  XNOR2_X1 prince_rounds_U197 ( .A(prince_rounds_SR_Inv_Result_s3[11]), .B(
        prince_rounds_n56), .ZN(prince_rounds_Output_s3[27]) );
  XNOR2_X1 prince_rounds_U196 ( .A(prince_rounds_SR_Inv_Result_s3[10]), .B(
        prince_rounds_n55), .ZN(prince_rounds_Output_s3[26]) );
  XNOR2_X1 prince_rounds_U195 ( .A(prince_rounds_SR_Inv_Result_s3[9]), .B(
        prince_rounds_n65), .ZN(prince_rounds_Output_s3[25]) );
  AOI22_X1 prince_rounds_U194 ( .A1(r[47]), .A2(prince_rounds_n49), .B1(r[63]), 
        .B2(prince_rounds_n48), .ZN(prince_rounds_n65) );
  XNOR2_X1 prince_rounds_U193 ( .A(prince_rounds_SR_Inv_Result_s3[8]), .B(
        prince_rounds_n64), .ZN(prince_rounds_Output_s3[24]) );
  AOI22_X1 prince_rounds_U192 ( .A1(r[46]), .A2(prince_rounds_n47), .B1(r[62]), 
        .B2(prince_rounds_n46), .ZN(prince_rounds_n64) );
  XNOR2_X1 prince_rounds_U191 ( .A(prince_rounds_SR_Inv_Result_s3[55]), .B(
        prince_rounds_n63), .ZN(prince_rounds_Output_s3[23]) );
  AOI22_X1 prince_rounds_U190 ( .A1(r[45]), .A2(prince_rounds_n45), .B1(r[61]), 
        .B2(prince_rounds_n44), .ZN(prince_rounds_n63) );
  XNOR2_X1 prince_rounds_U189 ( .A(prince_rounds_SR_Inv_Result_s3[54]), .B(
        prince_rounds_n62), .ZN(prince_rounds_Output_s3[22]) );
  AOI22_X1 prince_rounds_U188 ( .A1(r[44]), .A2(prince_rounds_n43), .B1(r[60]), 
        .B2(prince_rounds_n42), .ZN(prince_rounds_n62) );
  XNOR2_X1 prince_rounds_U187 ( .A(prince_rounds_SR_Inv_Result_s3[53]), .B(
        prince_rounds_n57), .ZN(prince_rounds_Output_s3[21]) );
  AOI22_X1 prince_rounds_U186 ( .A1(r[43]), .A2(prince_rounds_n41), .B1(r[59]), 
        .B2(prince_rounds_n40), .ZN(prince_rounds_n57) );
  XNOR2_X1 prince_rounds_U185 ( .A(prince_rounds_SR_Inv_Result_s3[52]), .B(
        prince_rounds_n54), .ZN(prince_rounds_Output_s3[20]) );
  AOI22_X1 prince_rounds_U184 ( .A1(r[42]), .A2(prince_rounds_n39), .B1(r[58]), 
        .B2(prince_rounds_n38), .ZN(prince_rounds_n54) );
  XNOR2_X1 prince_rounds_U183 ( .A(prince_rounds_SR_Inv_Result_s3[17]), .B(
        prince_rounds_n51), .ZN(prince_rounds_Output_s3[1]) );
  XNOR2_X1 prince_rounds_U182 ( .A(prince_rounds_SR_Inv_Result_s3[35]), .B(
        prince_rounds_n53), .ZN(prince_rounds_Output_s3[19]) );
  AOI22_X1 prince_rounds_U181 ( .A1(r[41]), .A2(prince_rounds_n37), .B1(r[57]), 
        .B2(prince_rounds_n36), .ZN(prince_rounds_n53) );
  XNOR2_X1 prince_rounds_U180 ( .A(prince_rounds_SR_Inv_Result_s3[34]), .B(
        prince_rounds_n52), .ZN(prince_rounds_Output_s3[18]) );
  AOI22_X1 prince_rounds_U179 ( .A1(r[40]), .A2(prince_rounds_n35), .B1(r[56]), 
        .B2(prince_rounds_n34), .ZN(prince_rounds_n52) );
  XNOR2_X1 prince_rounds_U178 ( .A(prince_rounds_SR_Inv_Result_s3[33]), .B(
        prince_rounds_n51), .ZN(prince_rounds_Output_s3[17]) );
  AOI22_X1 prince_rounds_U177 ( .A1(r[39]), .A2(prince_rounds_n33), .B1(r[55]), 
        .B2(prince_rounds_n32), .ZN(prince_rounds_n51) );
  XNOR2_X1 prince_rounds_U176 ( .A(prince_rounds_SR_Inv_Result_s3[32]), .B(
        prince_rounds_n50), .ZN(prince_rounds_Output_s3[16]) );
  XNOR2_X1 prince_rounds_U175 ( .A(prince_rounds_SR_Inv_Result_s3[15]), .B(
        prince_rounds_n61), .ZN(prince_rounds_Output_s3[15]) );
  AOI22_X1 prince_rounds_U174 ( .A1(r[53]), .A2(prince_rounds_n31), .B1(r[69]), 
        .B2(prince_rounds_n30), .ZN(prince_rounds_n61) );
  XNOR2_X1 prince_rounds_U173 ( .A(prince_rounds_SR_Inv_Result_s3[14]), .B(
        prince_rounds_n60), .ZN(prince_rounds_Output_s3[14]) );
  AOI22_X1 prince_rounds_U172 ( .A1(r[52]), .A2(prince_rounds_n29), .B1(r[68]), 
        .B2(prince_rounds_n28), .ZN(prince_rounds_n60) );
  XNOR2_X1 prince_rounds_U171 ( .A(prince_rounds_SR_Inv_Result_s3[13]), .B(
        prince_rounds_n59), .ZN(prince_rounds_Output_s3[13]) );
  AOI22_X1 prince_rounds_U170 ( .A1(r[51]), .A2(prince_rounds_n27), .B1(r[67]), 
        .B2(prince_rounds_n26), .ZN(prince_rounds_n59) );
  XNOR2_X1 prince_rounds_U169 ( .A(prince_rounds_SR_Inv_Result_s3[12]), .B(
        prince_rounds_n58), .ZN(prince_rounds_Output_s3[12]) );
  AOI22_X1 prince_rounds_U168 ( .A1(r[50]), .A2(prince_rounds_n25), .B1(r[66]), 
        .B2(prince_rounds_n24), .ZN(prince_rounds_n58) );
  XNOR2_X1 prince_rounds_U167 ( .A(prince_rounds_SR_Inv_Result_s3[59]), .B(
        prince_rounds_n56), .ZN(prince_rounds_Output_s3[11]) );
  AOI22_X1 prince_rounds_U166 ( .A1(r[49]), .A2(prince_rounds_n23), .B1(r[65]), 
        .B2(prince_rounds_n22), .ZN(prince_rounds_n56) );
  XNOR2_X1 prince_rounds_U165 ( .A(prince_rounds_SR_Inv_Result_s3[58]), .B(
        prince_rounds_n55), .ZN(prince_rounds_Output_s3[10]) );
  AOI22_X1 prince_rounds_U164 ( .A1(r[48]), .A2(prince_rounds_n21), .B1(r[64]), 
        .B2(prince_rounds_n20), .ZN(prince_rounds_n55) );
  XNOR2_X1 prince_rounds_U163 ( .A(prince_rounds_SR_Inv_Result_s3[16]), .B(
        prince_rounds_n50), .ZN(prince_rounds_Output_s3[0]) );
  AOI22_X1 prince_rounds_U162 ( .A1(r[38]), .A2(prince_rounds_n19), .B1(r[54]), 
        .B2(prince_rounds_n18), .ZN(prince_rounds_n50) );
  XNOR2_X1 prince_rounds_U161 ( .A(prince_rounds_SR_Inv_Result_s2[57]), .B(
        prince_rounds_n49), .ZN(prince_rounds_Output_s2[9]) );
  XNOR2_X1 prince_rounds_U160 ( .A(prince_rounds_SR_Inv_Result_s2[56]), .B(
        prince_rounds_n47), .ZN(prince_rounds_Output_s2[8]) );
  XNOR2_X1 prince_rounds_U159 ( .A(prince_rounds_SR_Inv_Result_s2[39]), .B(
        prince_rounds_n45), .ZN(prince_rounds_Output_s2[7]) );
  XNOR2_X1 prince_rounds_U158 ( .A(prince_rounds_SR_Inv_Result_s2[38]), .B(
        prince_rounds_n43), .ZN(prince_rounds_Output_s2[6]) );
  XNOR2_X1 prince_rounds_U157 ( .A(prince_rounds_SR_Inv_Result_s2[63]), .B(
        prince_rounds_n31), .ZN(prince_rounds_Output_s2[63]) );
  XNOR2_X1 prince_rounds_U156 ( .A(prince_rounds_SR_Inv_Result_s2[62]), .B(
        prince_rounds_n29), .ZN(prince_rounds_Output_s2[62]) );
  XNOR2_X1 prince_rounds_U155 ( .A(prince_rounds_SR_Inv_Result_s2[61]), .B(
        prince_rounds_n27), .ZN(prince_rounds_Output_s2[61]) );
  XNOR2_X1 prince_rounds_U154 ( .A(prince_rounds_SR_Inv_Result_s2[60]), .B(
        prince_rounds_n25), .ZN(prince_rounds_Output_s2[60]) );
  XNOR2_X1 prince_rounds_U153 ( .A(prince_rounds_SR_Inv_Result_s2[37]), .B(
        prince_rounds_n41), .ZN(prince_rounds_Output_s2[5]) );
  XNOR2_X1 prince_rounds_U152 ( .A(prince_rounds_SR_Inv_Result_s2[43]), .B(
        prince_rounds_n23), .ZN(prince_rounds_Output_s2[59]) );
  XNOR2_X1 prince_rounds_U151 ( .A(prince_rounds_SR_Inv_Result_s2[42]), .B(
        prince_rounds_n21), .ZN(prince_rounds_Output_s2[58]) );
  XNOR2_X1 prince_rounds_U150 ( .A(prince_rounds_SR_Inv_Result_s2[41]), .B(
        prince_rounds_n49), .ZN(prince_rounds_Output_s2[57]) );
  XNOR2_X1 prince_rounds_U149 ( .A(prince_rounds_SR_Inv_Result_s2[40]), .B(
        prince_rounds_n47), .ZN(prince_rounds_Output_s2[56]) );
  XNOR2_X1 prince_rounds_U148 ( .A(prince_rounds_SR_Inv_Result_s2[23]), .B(
        prince_rounds_n45), .ZN(prince_rounds_Output_s2[55]) );
  XNOR2_X1 prince_rounds_U147 ( .A(prince_rounds_SR_Inv_Result_s2[22]), .B(
        prince_rounds_n43), .ZN(prince_rounds_Output_s2[54]) );
  XNOR2_X1 prince_rounds_U146 ( .A(prince_rounds_SR_Inv_Result_s2[21]), .B(
        prince_rounds_n41), .ZN(prince_rounds_Output_s2[53]) );
  XNOR2_X1 prince_rounds_U145 ( .A(prince_rounds_SR_Inv_Result_s2[20]), .B(
        prince_rounds_n39), .ZN(prince_rounds_Output_s2[52]) );
  XNOR2_X1 prince_rounds_U144 ( .A(prince_rounds_SR_Inv_Result_s2[3]), .B(
        prince_rounds_n37), .ZN(prince_rounds_Output_s2[51]) );
  XNOR2_X1 prince_rounds_U143 ( .A(prince_rounds_SR_Inv_Result_s2[2]), .B(
        prince_rounds_n35), .ZN(prince_rounds_Output_s2[50]) );
  XNOR2_X1 prince_rounds_U142 ( .A(prince_rounds_SR_Inv_Result_s2[36]), .B(
        prince_rounds_n39), .ZN(prince_rounds_Output_s2[4]) );
  XNOR2_X1 prince_rounds_U141 ( .A(prince_rounds_SR_Inv_Result_s2[1]), .B(
        prince_rounds_n33), .ZN(prince_rounds_Output_s2[49]) );
  XNOR2_X1 prince_rounds_U140 ( .A(prince_rounds_SR_Inv_Result_s2[0]), .B(
        prince_rounds_n19), .ZN(prince_rounds_Output_s2[48]) );
  XNOR2_X1 prince_rounds_U139 ( .A(prince_rounds_SR_Inv_Result_s2[47]), .B(
        prince_rounds_n31), .ZN(prince_rounds_Output_s2[47]) );
  XNOR2_X1 prince_rounds_U138 ( .A(prince_rounds_SR_Inv_Result_s2[46]), .B(
        prince_rounds_n29), .ZN(prince_rounds_Output_s2[46]) );
  XNOR2_X1 prince_rounds_U137 ( .A(prince_rounds_SR_Inv_Result_s2[45]), .B(
        prince_rounds_n27), .ZN(prince_rounds_Output_s2[45]) );
  XNOR2_X1 prince_rounds_U136 ( .A(prince_rounds_SR_Inv_Result_s2[44]), .B(
        prince_rounds_n25), .ZN(prince_rounds_Output_s2[44]) );
  XNOR2_X1 prince_rounds_U135 ( .A(prince_rounds_SR_Inv_Result_s2[27]), .B(
        prince_rounds_n23), .ZN(prince_rounds_Output_s2[43]) );
  XNOR2_X1 prince_rounds_U134 ( .A(prince_rounds_SR_Inv_Result_s2[26]), .B(
        prince_rounds_n21), .ZN(prince_rounds_Output_s2[42]) );
  XNOR2_X1 prince_rounds_U133 ( .A(prince_rounds_SR_Inv_Result_s2[25]), .B(
        prince_rounds_n49), .ZN(prince_rounds_Output_s2[41]) );
  XNOR2_X1 prince_rounds_U132 ( .A(prince_rounds_SR_Inv_Result_s2[24]), .B(
        prince_rounds_n47), .ZN(prince_rounds_Output_s2[40]) );
  XNOR2_X1 prince_rounds_U131 ( .A(prince_rounds_SR_Inv_Result_s2[19]), .B(
        prince_rounds_n37), .ZN(prince_rounds_Output_s2[3]) );
  XNOR2_X1 prince_rounds_U130 ( .A(prince_rounds_SR_Inv_Result_s2[7]), .B(
        prince_rounds_n45), .ZN(prince_rounds_Output_s2[39]) );
  XNOR2_X1 prince_rounds_U129 ( .A(prince_rounds_SR_Inv_Result_s2[6]), .B(
        prince_rounds_n43), .ZN(prince_rounds_Output_s2[38]) );
  XNOR2_X1 prince_rounds_U128 ( .A(prince_rounds_SR_Inv_Result_s2[5]), .B(
        prince_rounds_n41), .ZN(prince_rounds_Output_s2[37]) );
  XNOR2_X1 prince_rounds_U127 ( .A(prince_rounds_SR_Inv_Result_s2[4]), .B(
        prince_rounds_n39), .ZN(prince_rounds_Output_s2[36]) );
  XNOR2_X1 prince_rounds_U126 ( .A(prince_rounds_SR_Inv_Result_s2[51]), .B(
        prince_rounds_n37), .ZN(prince_rounds_Output_s2[35]) );
  XNOR2_X1 prince_rounds_U125 ( .A(prince_rounds_SR_Inv_Result_s2[50]), .B(
        prince_rounds_n35), .ZN(prince_rounds_Output_s2[34]) );
  XNOR2_X1 prince_rounds_U124 ( .A(prince_rounds_SR_Inv_Result_s2[49]), .B(
        prince_rounds_n33), .ZN(prince_rounds_Output_s2[33]) );
  XNOR2_X1 prince_rounds_U123 ( .A(prince_rounds_SR_Inv_Result_s2[48]), .B(
        prince_rounds_n19), .ZN(prince_rounds_Output_s2[32]) );
  XNOR2_X1 prince_rounds_U122 ( .A(prince_rounds_SR_Inv_Result_s2[31]), .B(
        prince_rounds_n31), .ZN(prince_rounds_Output_s2[31]) );
  XNOR2_X1 prince_rounds_U121 ( .A(prince_rounds_SR_Inv_Result_s2[30]), .B(
        prince_rounds_n29), .ZN(prince_rounds_Output_s2[30]) );
  XNOR2_X1 prince_rounds_U120 ( .A(prince_rounds_SR_Inv_Result_s2[18]), .B(
        prince_rounds_n35), .ZN(prince_rounds_Output_s2[2]) );
  XNOR2_X1 prince_rounds_U119 ( .A(prince_rounds_SR_Inv_Result_s2[29]), .B(
        prince_rounds_n27), .ZN(prince_rounds_Output_s2[29]) );
  XNOR2_X1 prince_rounds_U118 ( .A(prince_rounds_SR_Inv_Result_s2[28]), .B(
        prince_rounds_n25), .ZN(prince_rounds_Output_s2[28]) );
  XNOR2_X1 prince_rounds_U117 ( .A(prince_rounds_SR_Inv_Result_s2[11]), .B(
        prince_rounds_n23), .ZN(prince_rounds_Output_s2[27]) );
  XNOR2_X1 prince_rounds_U116 ( .A(prince_rounds_SR_Inv_Result_s2[10]), .B(
        prince_rounds_n21), .ZN(prince_rounds_Output_s2[26]) );
  XNOR2_X1 prince_rounds_U115 ( .A(prince_rounds_SR_Inv_Result_s2[9]), .B(
        prince_rounds_n49), .ZN(prince_rounds_Output_s2[25]) );
  XNOR2_X1 prince_rounds_U114 ( .A(prince_rounds_SR_Inv_Result_s2[8]), .B(
        prince_rounds_n47), .ZN(prince_rounds_Output_s2[24]) );
  XNOR2_X1 prince_rounds_U113 ( .A(prince_rounds_SR_Inv_Result_s2[55]), .B(
        prince_rounds_n45), .ZN(prince_rounds_Output_s2[23]) );
  XNOR2_X1 prince_rounds_U112 ( .A(prince_rounds_SR_Inv_Result_s2[54]), .B(
        prince_rounds_n43), .ZN(prince_rounds_Output_s2[22]) );
  XNOR2_X1 prince_rounds_U111 ( .A(prince_rounds_SR_Inv_Result_s2[53]), .B(
        prince_rounds_n41), .ZN(prince_rounds_Output_s2[21]) );
  XNOR2_X1 prince_rounds_U110 ( .A(prince_rounds_SR_Inv_Result_s2[52]), .B(
        prince_rounds_n39), .ZN(prince_rounds_Output_s2[20]) );
  XNOR2_X1 prince_rounds_U109 ( .A(prince_rounds_SR_Inv_Result_s2[17]), .B(
        prince_rounds_n33), .ZN(prince_rounds_Output_s2[1]) );
  XNOR2_X1 prince_rounds_U108 ( .A(prince_rounds_SR_Inv_Result_s2[35]), .B(
        prince_rounds_n37), .ZN(prince_rounds_Output_s2[19]) );
  XNOR2_X1 prince_rounds_U107 ( .A(prince_rounds_SR_Inv_Result_s2[34]), .B(
        prince_rounds_n35), .ZN(prince_rounds_Output_s2[18]) );
  XNOR2_X1 prince_rounds_U106 ( .A(prince_rounds_SR_Inv_Result_s2[33]), .B(
        prince_rounds_n33), .ZN(prince_rounds_Output_s2[17]) );
  XNOR2_X1 prince_rounds_U105 ( .A(prince_rounds_SR_Inv_Result_s2[32]), .B(
        prince_rounds_n19), .ZN(prince_rounds_Output_s2[16]) );
  XNOR2_X1 prince_rounds_U104 ( .A(prince_rounds_SR_Inv_Result_s2[15]), .B(
        prince_rounds_n31), .ZN(prince_rounds_Output_s2[15]) );
  XNOR2_X1 prince_rounds_U103 ( .A(prince_rounds_SR_Inv_Result_s2[14]), .B(
        prince_rounds_n29), .ZN(prince_rounds_Output_s2[14]) );
  XNOR2_X1 prince_rounds_U102 ( .A(prince_rounds_SR_Inv_Result_s2[13]), .B(
        prince_rounds_n27), .ZN(prince_rounds_Output_s2[13]) );
  XNOR2_X1 prince_rounds_U101 ( .A(prince_rounds_SR_Inv_Result_s2[12]), .B(
        prince_rounds_n25), .ZN(prince_rounds_Output_s2[12]) );
  XNOR2_X1 prince_rounds_U100 ( .A(prince_rounds_SR_Inv_Result_s2[59]), .B(
        prince_rounds_n23), .ZN(prince_rounds_Output_s2[11]) );
  XNOR2_X1 prince_rounds_U99 ( .A(prince_rounds_SR_Inv_Result_s2[58]), .B(
        prince_rounds_n21), .ZN(prince_rounds_Output_s2[10]) );
  XNOR2_X1 prince_rounds_U98 ( .A(prince_rounds_SR_Inv_Result_s2[16]), .B(
        prince_rounds_n19), .ZN(prince_rounds_Output_s2[0]) );
  XNOR2_X1 prince_rounds_U97 ( .A(prince_rounds_SR_Inv_Result_s1[57]), .B(
        prince_rounds_n48), .ZN(prince_rounds_Output_s1[9]) );
  XNOR2_X1 prince_rounds_U96 ( .A(prince_rounds_SR_Inv_Result_s1[56]), .B(
        prince_rounds_n46), .ZN(prince_rounds_Output_s1[8]) );
  XNOR2_X1 prince_rounds_U95 ( .A(prince_rounds_SR_Inv_Result_s1[39]), .B(
        prince_rounds_n44), .ZN(prince_rounds_Output_s1[7]) );
  XNOR2_X1 prince_rounds_U94 ( .A(prince_rounds_SR_Inv_Result_s1[38]), .B(
        prince_rounds_n42), .ZN(prince_rounds_Output_s1[6]) );
  XNOR2_X1 prince_rounds_U93 ( .A(prince_rounds_SR_Inv_Result_s1[63]), .B(
        prince_rounds_n30), .ZN(prince_rounds_Output_s1[63]) );
  XNOR2_X1 prince_rounds_U92 ( .A(prince_rounds_SR_Inv_Result_s1[62]), .B(
        prince_rounds_n28), .ZN(prince_rounds_Output_s1[62]) );
  XNOR2_X1 prince_rounds_U91 ( .A(prince_rounds_SR_Inv_Result_s1[61]), .B(
        prince_rounds_n26), .ZN(prince_rounds_Output_s1[61]) );
  XNOR2_X1 prince_rounds_U90 ( .A(prince_rounds_SR_Inv_Result_s1[60]), .B(
        prince_rounds_n24), .ZN(prince_rounds_Output_s1[60]) );
  XNOR2_X1 prince_rounds_U89 ( .A(prince_rounds_SR_Inv_Result_s1[37]), .B(
        prince_rounds_n40), .ZN(prince_rounds_Output_s1[5]) );
  XNOR2_X1 prince_rounds_U88 ( .A(prince_rounds_SR_Inv_Result_s1[43]), .B(
        prince_rounds_n22), .ZN(prince_rounds_Output_s1[59]) );
  XNOR2_X1 prince_rounds_U87 ( .A(prince_rounds_SR_Inv_Result_s1[42]), .B(
        prince_rounds_n20), .ZN(prince_rounds_Output_s1[58]) );
  XNOR2_X1 prince_rounds_U86 ( .A(prince_rounds_SR_Inv_Result_s1[41]), .B(
        prince_rounds_n48), .ZN(prince_rounds_Output_s1[57]) );
  XNOR2_X1 prince_rounds_U85 ( .A(prince_rounds_SR_Inv_Result_s1[40]), .B(
        prince_rounds_n46), .ZN(prince_rounds_Output_s1[56]) );
  XNOR2_X1 prince_rounds_U84 ( .A(prince_rounds_SR_Inv_Result_s1[23]), .B(
        prince_rounds_n44), .ZN(prince_rounds_Output_s1[55]) );
  XNOR2_X1 prince_rounds_U83 ( .A(prince_rounds_SR_Inv_Result_s1[22]), .B(
        prince_rounds_n42), .ZN(prince_rounds_Output_s1[54]) );
  XNOR2_X1 prince_rounds_U82 ( .A(prince_rounds_SR_Inv_Result_s1[21]), .B(
        prince_rounds_n40), .ZN(prince_rounds_Output_s1[53]) );
  XNOR2_X1 prince_rounds_U81 ( .A(prince_rounds_SR_Inv_Result_s1[20]), .B(
        prince_rounds_n38), .ZN(prince_rounds_Output_s1[52]) );
  XNOR2_X1 prince_rounds_U80 ( .A(prince_rounds_SR_Inv_Result_s1[3]), .B(
        prince_rounds_n36), .ZN(prince_rounds_Output_s1[51]) );
  XNOR2_X1 prince_rounds_U79 ( .A(prince_rounds_SR_Inv_Result_s1[2]), .B(
        prince_rounds_n34), .ZN(prince_rounds_Output_s1[50]) );
  XNOR2_X1 prince_rounds_U78 ( .A(prince_rounds_SR_Inv_Result_s1[36]), .B(
        prince_rounds_n38), .ZN(prince_rounds_Output_s1[4]) );
  XNOR2_X1 prince_rounds_U77 ( .A(prince_rounds_SR_Inv_Result_s1[1]), .B(
        prince_rounds_n32), .ZN(prince_rounds_Output_s1[49]) );
  XNOR2_X1 prince_rounds_U76 ( .A(prince_rounds_SR_Inv_Result_s1[0]), .B(
        prince_rounds_n18), .ZN(prince_rounds_Output_s1[48]) );
  XNOR2_X1 prince_rounds_U75 ( .A(prince_rounds_SR_Inv_Result_s1[47]), .B(
        prince_rounds_n30), .ZN(prince_rounds_Output_s1[47]) );
  XNOR2_X1 prince_rounds_U74 ( .A(prince_rounds_SR_Inv_Result_s1[46]), .B(
        prince_rounds_n28), .ZN(prince_rounds_Output_s1[46]) );
  XNOR2_X1 prince_rounds_U73 ( .A(prince_rounds_SR_Inv_Result_s1[45]), .B(
        prince_rounds_n26), .ZN(prince_rounds_Output_s1[45]) );
  XNOR2_X1 prince_rounds_U72 ( .A(prince_rounds_SR_Inv_Result_s1[44]), .B(
        prince_rounds_n24), .ZN(prince_rounds_Output_s1[44]) );
  XNOR2_X1 prince_rounds_U71 ( .A(prince_rounds_SR_Inv_Result_s1[27]), .B(
        prince_rounds_n22), .ZN(prince_rounds_Output_s1[43]) );
  XNOR2_X1 prince_rounds_U70 ( .A(prince_rounds_SR_Inv_Result_s1[26]), .B(
        prince_rounds_n20), .ZN(prince_rounds_Output_s1[42]) );
  XNOR2_X1 prince_rounds_U69 ( .A(prince_rounds_SR_Inv_Result_s1[25]), .B(
        prince_rounds_n48), .ZN(prince_rounds_Output_s1[41]) );
  XNOR2_X1 prince_rounds_U68 ( .A(prince_rounds_SR_Inv_Result_s1[24]), .B(
        prince_rounds_n46), .ZN(prince_rounds_Output_s1[40]) );
  XNOR2_X1 prince_rounds_U67 ( .A(prince_rounds_SR_Inv_Result_s1[19]), .B(
        prince_rounds_n36), .ZN(prince_rounds_Output_s1[3]) );
  XNOR2_X1 prince_rounds_U66 ( .A(prince_rounds_SR_Inv_Result_s1[7]), .B(
        prince_rounds_n44), .ZN(prince_rounds_Output_s1[39]) );
  XNOR2_X1 prince_rounds_U65 ( .A(prince_rounds_SR_Inv_Result_s1[6]), .B(
        prince_rounds_n42), .ZN(prince_rounds_Output_s1[38]) );
  XNOR2_X1 prince_rounds_U64 ( .A(prince_rounds_SR_Inv_Result_s1[5]), .B(
        prince_rounds_n40), .ZN(prince_rounds_Output_s1[37]) );
  XNOR2_X1 prince_rounds_U63 ( .A(prince_rounds_SR_Inv_Result_s1[4]), .B(
        prince_rounds_n38), .ZN(prince_rounds_Output_s1[36]) );
  XNOR2_X1 prince_rounds_U62 ( .A(prince_rounds_SR_Inv_Result_s1[51]), .B(
        prince_rounds_n36), .ZN(prince_rounds_Output_s1[35]) );
  XNOR2_X1 prince_rounds_U61 ( .A(prince_rounds_SR_Inv_Result_s1[50]), .B(
        prince_rounds_n34), .ZN(prince_rounds_Output_s1[34]) );
  XNOR2_X1 prince_rounds_U60 ( .A(prince_rounds_SR_Inv_Result_s1[49]), .B(
        prince_rounds_n32), .ZN(prince_rounds_Output_s1[33]) );
  XNOR2_X1 prince_rounds_U59 ( .A(prince_rounds_SR_Inv_Result_s1[48]), .B(
        prince_rounds_n18), .ZN(prince_rounds_Output_s1[32]) );
  XNOR2_X1 prince_rounds_U58 ( .A(prince_rounds_SR_Inv_Result_s1[31]), .B(
        prince_rounds_n30), .ZN(prince_rounds_Output_s1[31]) );
  XNOR2_X1 prince_rounds_U57 ( .A(prince_rounds_SR_Inv_Result_s1[30]), .B(
        prince_rounds_n28), .ZN(prince_rounds_Output_s1[30]) );
  XNOR2_X1 prince_rounds_U56 ( .A(prince_rounds_SR_Inv_Result_s1[18]), .B(
        prince_rounds_n34), .ZN(prince_rounds_Output_s1[2]) );
  XNOR2_X1 prince_rounds_U55 ( .A(prince_rounds_SR_Inv_Result_s1[29]), .B(
        prince_rounds_n26), .ZN(prince_rounds_Output_s1[29]) );
  XNOR2_X1 prince_rounds_U54 ( .A(prince_rounds_SR_Inv_Result_s1[28]), .B(
        prince_rounds_n24), .ZN(prince_rounds_Output_s1[28]) );
  XNOR2_X1 prince_rounds_U53 ( .A(prince_rounds_SR_Inv_Result_s1[11]), .B(
        prince_rounds_n22), .ZN(prince_rounds_Output_s1[27]) );
  XNOR2_X1 prince_rounds_U52 ( .A(prince_rounds_SR_Inv_Result_s1[10]), .B(
        prince_rounds_n20), .ZN(prince_rounds_Output_s1[26]) );
  XNOR2_X1 prince_rounds_U51 ( .A(prince_rounds_SR_Inv_Result_s1[9]), .B(
        prince_rounds_n48), .ZN(prince_rounds_Output_s1[25]) );
  XNOR2_X1 prince_rounds_U50 ( .A(prince_rounds_SR_Inv_Result_s1[8]), .B(
        prince_rounds_n46), .ZN(prince_rounds_Output_s1[24]) );
  XNOR2_X1 prince_rounds_U49 ( .A(prince_rounds_SR_Inv_Result_s1[55]), .B(
        prince_rounds_n44), .ZN(prince_rounds_Output_s1[23]) );
  XNOR2_X1 prince_rounds_U48 ( .A(prince_rounds_SR_Inv_Result_s1[54]), .B(
        prince_rounds_n42), .ZN(prince_rounds_Output_s1[22]) );
  XNOR2_X1 prince_rounds_U47 ( .A(prince_rounds_SR_Inv_Result_s1[53]), .B(
        prince_rounds_n40), .ZN(prince_rounds_Output_s1[21]) );
  XNOR2_X1 prince_rounds_U46 ( .A(prince_rounds_SR_Inv_Result_s1[52]), .B(
        prince_rounds_n38), .ZN(prince_rounds_Output_s1[20]) );
  XNOR2_X1 prince_rounds_U45 ( .A(prince_rounds_SR_Inv_Result_s1[17]), .B(
        prince_rounds_n32), .ZN(prince_rounds_Output_s1[1]) );
  XNOR2_X1 prince_rounds_U44 ( .A(prince_rounds_SR_Inv_Result_s1[35]), .B(
        prince_rounds_n36), .ZN(prince_rounds_Output_s1[19]) );
  XNOR2_X1 prince_rounds_U43 ( .A(prince_rounds_SR_Inv_Result_s1[34]), .B(
        prince_rounds_n34), .ZN(prince_rounds_Output_s1[18]) );
  XNOR2_X1 prince_rounds_U42 ( .A(prince_rounds_SR_Inv_Result_s1[33]), .B(
        prince_rounds_n32), .ZN(prince_rounds_Output_s1[17]) );
  XNOR2_X1 prince_rounds_U41 ( .A(prince_rounds_SR_Inv_Result_s1[32]), .B(
        prince_rounds_n18), .ZN(prince_rounds_Output_s1[16]) );
  XNOR2_X1 prince_rounds_U40 ( .A(prince_rounds_SR_Inv_Result_s1[15]), .B(
        prince_rounds_n30), .ZN(prince_rounds_Output_s1[15]) );
  XNOR2_X1 prince_rounds_U39 ( .A(prince_rounds_SR_Inv_Result_s1[14]), .B(
        prince_rounds_n28), .ZN(prince_rounds_Output_s1[14]) );
  XNOR2_X1 prince_rounds_U38 ( .A(prince_rounds_SR_Inv_Result_s1[13]), .B(
        prince_rounds_n26), .ZN(prince_rounds_Output_s1[13]) );
  XNOR2_X1 prince_rounds_U37 ( .A(prince_rounds_SR_Inv_Result_s1[12]), .B(
        prince_rounds_n24), .ZN(prince_rounds_Output_s1[12]) );
  XNOR2_X1 prince_rounds_U36 ( .A(prince_rounds_SR_Inv_Result_s1[59]), .B(
        prince_rounds_n22), .ZN(prince_rounds_Output_s1[11]) );
  XNOR2_X1 prince_rounds_U35 ( .A(prince_rounds_SR_Inv_Result_s1[58]), .B(
        prince_rounds_n20), .ZN(prince_rounds_Output_s1[10]) );
  XNOR2_X1 prince_rounds_U34 ( .A(prince_rounds_SR_Inv_Result_s1[16]), .B(
        prince_rounds_n18), .ZN(prince_rounds_Output_s1[0]) );
  INV_X1 prince_rounds_U33 ( .A(r[45]), .ZN(prince_rounds_n44) );
  INV_X1 prince_rounds_U32 ( .A(r[54]), .ZN(prince_rounds_n19) );
  INV_X1 prince_rounds_U31 ( .A(r[41]), .ZN(prince_rounds_n36) );
  INV_X1 prince_rounds_U30 ( .A(r[40]), .ZN(prince_rounds_n34) );
  INV_X1 prince_rounds_U29 ( .A(r[63]), .ZN(prince_rounds_n49) );
  INV_X1 prince_rounds_U28 ( .A(r[62]), .ZN(prince_rounds_n47) );
  INV_X1 prince_rounds_U27 ( .A(r[58]), .ZN(prince_rounds_n39) );
  INV_X1 prince_rounds_U26 ( .A(r[65]), .ZN(prince_rounds_n23) );
  INV_X1 prince_rounds_U25 ( .A(r[66]), .ZN(prince_rounds_n25) );
  INV_X1 prince_rounds_U24 ( .A(r[60]), .ZN(prince_rounds_n43) );
  INV_X1 prince_rounds_U23 ( .A(r[46]), .ZN(prince_rounds_n46) );
  INV_X1 prince_rounds_U22 ( .A(r[50]), .ZN(prince_rounds_n24) );
  INV_X1 prince_rounds_U21 ( .A(r[47]), .ZN(prince_rounds_n48) );
  INV_X1 prince_rounds_U20 ( .A(r[67]), .ZN(prince_rounds_n27) );
  INV_X1 prince_rounds_U19 ( .A(r[68]), .ZN(prince_rounds_n29) );
  INV_X1 prince_rounds_U18 ( .A(r[64]), .ZN(prince_rounds_n21) );
  INV_X1 prince_rounds_U17 ( .A(r[55]), .ZN(prince_rounds_n33) );
  INV_X1 prince_rounds_U16 ( .A(r[69]), .ZN(prince_rounds_n31) );
  INV_X1 prince_rounds_U15 ( .A(r[56]), .ZN(prince_rounds_n35) );
  INV_X1 prince_rounds_U14 ( .A(r[57]), .ZN(prince_rounds_n37) );
  INV_X1 prince_rounds_U13 ( .A(r[39]), .ZN(prince_rounds_n32) );
  INV_X1 prince_rounds_U12 ( .A(r[59]), .ZN(prince_rounds_n41) );
  INV_X1 prince_rounds_U11 ( .A(r[38]), .ZN(prince_rounds_n18) );
  INV_X1 prince_rounds_U10 ( .A(r[61]), .ZN(prince_rounds_n45) );
  INV_X1 prince_rounds_U9 ( .A(r[53]), .ZN(prince_rounds_n30) );
  INV_X1 prince_rounds_U8 ( .A(r[52]), .ZN(prince_rounds_n28) );
  INV_X1 prince_rounds_U7 ( .A(r[51]), .ZN(prince_rounds_n26) );
  INV_X1 prince_rounds_U6 ( .A(r[48]), .ZN(prince_rounds_n20) );
  INV_X1 prince_rounds_U5 ( .A(r[49]), .ZN(prince_rounds_n22) );
  INV_X1 prince_rounds_U4 ( .A(r[43]), .ZN(prince_rounds_n40) );
  INV_X1 prince_rounds_U3 ( .A(r[44]), .ZN(prince_rounds_n42) );
  INV_X1 prince_rounds_U2 ( .A(r[42]), .ZN(prince_rounds_n38) );
  NAND2_X1 prince_rounds_constant_MUX_U87 ( .A1(prince_rounds_constant_MUX_n46), .A2(prince_rounds_constant_MUX_n45), .ZN(prince_rounds_round_Constant[8]) );
  NAND2_X1 prince_rounds_constant_MUX_U86 ( .A1(prince_rounds_constant_MUX_n44), .A2(prince_rounds_constant_MUX_n43), .ZN(prince_rounds_round_Constant[18])
         );
  NAND4_X1 prince_rounds_constant_MUX_U85 ( .A1(prince_rounds_constant_MUX_n42), .A2(prince_rounds_constant_MUX_n41), .A3(prince_rounds_constant_MUX_n40), 
        .A4(prince_rounds_constant_MUX_n39), .ZN(
        prince_rounds_round_Constant[33]) );
  NAND4_X1 prince_rounds_constant_MUX_U84 ( .A1(prince_rounds_constant_MUX_n38), .A2(prince_rounds_constant_MUX_n37), .A3(prince_rounds_constant_MUX_n40), 
        .A4(prince_rounds_constant_MUX_n39), .ZN(
        prince_rounds_round_Constant[4]) );
  NAND2_X1 prince_rounds_constant_MUX_U83 ( .A1(prince_rounds_constant_MUX_n36), .A2(prince_rounds_constant_MUX_n35), .ZN(prince_rounds_round_Constant[50])
         );
  NAND2_X1 prince_rounds_constant_MUX_U82 ( .A1(prince_rounds_constant_MUX_n34), .A2(prince_rounds_constant_MUX_n40), .ZN(prince_rounds_round_Constant[34])
         );
  NAND3_X1 prince_rounds_constant_MUX_U81 ( .A1(prince_rounds_constant_MUX_n33), .A2(prince_rounds_constant_MUX_n32), .A3(prince_rounds_constant_MUX_n43), 
        .ZN(prince_rounds_round_Constant[14]) );
  OR2_X1 prince_rounds_constant_MUX_U80 ( .A1(prince_rounds_round_Constant[49]), .A2(prince_rounds_round_Constant[48]), .ZN(prince_rounds_round_Constant[13])
         );
  NAND2_X1 prince_rounds_constant_MUX_U79 ( .A1(prince_rounds_constant_MUX_n31), .A2(prince_rounds_constant_MUX_n40), .ZN(prince_rounds_round_Constant[37])
         );
  NAND2_X1 prince_rounds_constant_MUX_U78 ( .A1(prince_rounds_constant_MUX_n38), .A2(prince_rounds_constant_MUX_n35), .ZN(prince_rounds_round_Constant[53])
         );
  NAND4_X1 prince_rounds_constant_MUX_U77 ( .A1(prince_rounds_constant_MUX_n36), .A2(prince_rounds_constant_MUX_n37), .A3(prince_rounds_constant_MUX_n40), 
        .A4(prince_rounds_constant_MUX_n39), .ZN(
        prince_rounds_round_Constant[63]) );
  NAND2_X1 prince_rounds_constant_MUX_U76 ( .A1(prince_rounds_constant_MUX_n38), .A2(prince_rounds_constant_MUX_n30), .ZN(prince_rounds_round_Constant[62])
         );
  NAND2_X1 prince_rounds_constant_MUX_U75 ( .A1(prince_rounds_constant_MUX_n29), .A2(prince_rounds_constant_MUX_n46), .ZN(prince_rounds_round_Constant[61])
         );
  NAND2_X1 prince_rounds_constant_MUX_U74 ( .A1(prince_rounds_constant_MUX_n46), .A2(prince_rounds_constant_MUX_n28), .ZN(prince_rounds_round_Constant[58])
         );
  INV_X1 prince_rounds_constant_MUX_U73 ( .A(prince_rounds_round_Constant[38]), 
        .ZN(prince_rounds_constant_MUX_n28) );
  NAND2_X1 prince_rounds_constant_MUX_U72 ( .A1(prince_rounds_constant_MUX_n27), .A2(prince_rounds_constant_MUX_n37), .ZN(prince_rounds_round_Constant[55])
         );
  NAND2_X1 prince_rounds_constant_MUX_U71 ( .A1(prince_rounds_constant_MUX_n31), .A2(prince_rounds_constant_MUX_n32), .ZN(prince_rounds_round_Constant[51])
         );
  NOR2_X1 prince_rounds_constant_MUX_U70 ( .A1(prince_rounds_constant_MUX_n26), 
        .A2(prince_rounds_constant_MUX_n25), .ZN(
        prince_rounds_constant_MUX_n31) );
  NAND3_X1 prince_rounds_constant_MUX_U69 ( .A1(prince_rounds_constant_MUX_n42), .A2(prince_rounds_constant_MUX_n39), .A3(prince_rounds_constant_MUX_n24), 
        .ZN(prince_rounds_constant_MUX_n25) );
  NAND2_X1 prince_rounds_constant_MUX_U68 ( .A1(prince_rounds_constant_MUX_n23), .A2(prince_rounds_constant_MUX_n46), .ZN(prince_rounds_round_Constant[48])
         );
  NAND2_X1 prince_rounds_constant_MUX_U67 ( .A1(prince_rounds_constant_MUX_n22), .A2(prince_rounds_constant_MUX_n23), .ZN(prince_rounds_round_Constant[47])
         );
  NAND2_X1 prince_rounds_constant_MUX_U66 ( .A1(prince_rounds_constant_MUX_n41), .A2(prince_rounds_constant_MUX_n44), .ZN(prince_rounds_round_Constant[45])
         );
  NAND2_X1 prince_rounds_constant_MUX_U65 ( .A1(prince_rounds_constant_MUX_n22), .A2(prince_rounds_constant_MUX_n46), .ZN(prince_rounds_round_Constant[44])
         );
  NAND2_X1 prince_rounds_constant_MUX_U64 ( .A1(prince_rounds_constant_MUX_n20), .A2(prince_rounds_constant_MUX_n19), .ZN(prince_rounds_constant_MUX_n39) );
  NAND2_X1 prince_rounds_constant_MUX_U63 ( .A1(prince_rounds_constant_MUX_n18), .A2(prince_rounds_constant_MUX_n32), .ZN(prince_rounds_round_Constant[43])
         );
  OR2_X1 prince_rounds_constant_MUX_U62 ( .A1(prince_rounds_round_Constant[49]), .A2(prince_rounds_round_Constant[60]), .ZN(prince_rounds_round_Constant[41])
         );
  NAND2_X1 prince_rounds_constant_MUX_U61 ( .A1(prince_rounds_constant_MUX_n23), .A2(prince_rounds_constant_MUX_n29), .ZN(prince_rounds_round_Constant[60])
         );
  NAND2_X1 prince_rounds_constant_MUX_U60 ( .A1(prince_rounds_constant_MUX_n22), .A2(prince_rounds_constant_MUX_n29), .ZN(prince_rounds_round_Constant[59])
         );
  INV_X1 prince_rounds_constant_MUX_U59 ( .A(prince_rounds_round_Constant[54]), 
        .ZN(prince_rounds_constant_MUX_n29) );
  INV_X1 prince_rounds_constant_MUX_U58 ( .A(prince_rounds_round_Constant[49]), 
        .ZN(prince_rounds_constant_MUX_n22) );
  NAND2_X1 prince_rounds_constant_MUX_U57 ( .A1(prince_rounds_constant_MUX_n32), .A2(prince_rounds_constant_MUX_n40), .ZN(prince_rounds_round_Constant[49])
         );
  NAND2_X1 prince_rounds_constant_MUX_U56 ( .A1(prince_rounds_constant_MUX_n35), .A2(prince_rounds_constant_MUX_n41), .ZN(prince_rounds_round_Constant[39])
         );
  NAND2_X1 prince_rounds_constant_MUX_U55 ( .A1(prince_rounds_constant_MUX_n35), .A2(prince_rounds_constant_MUX_n43), .ZN(prince_rounds_round_Constant[36])
         );
  AND3_X1 prince_rounds_constant_MUX_U54 ( .A1(prince_rounds_constant_MUX_n32), 
        .A2(prince_rounds_constant_MUX_n21), .A3(
        prince_rounds_constant_MUX_n37), .ZN(prince_rounds_constant_MUX_n35)
         );
  INV_X1 prince_rounds_constant_MUX_U53 ( .A(prince_rounds_constant_MUX_n17), 
        .ZN(prince_rounds_constant_MUX_n37) );
  NAND2_X1 prince_rounds_constant_MUX_U52 ( .A1(prince_rounds_constant_MUX_n36), .A2(prince_rounds_constant_MUX_n30), .ZN(prince_rounds_round_Constant[32])
         );
  AOI21_X1 prince_rounds_constant_MUX_U51 ( .B1(prince_rounds_constant_MUX_n16), .B2(prince_rounds_constant_MUX_n15), .A(prince_rounds_constant_MUX_n17), 
        .ZN(prince_rounds_constant_MUX_n30) );
  NAND2_X1 prince_rounds_constant_MUX_U50 ( .A1(prince_rounds_constant_MUX_n14), .A2(prince_rounds_constant_MUX_n27), .ZN(prince_rounds_round_Constant[29])
         );
  NAND2_X1 prince_rounds_constant_MUX_U49 ( .A1(prince_rounds_constant_MUX_n38), .A2(prince_rounds_constant_MUX_n44), .ZN(prince_rounds_round_Constant[27])
         );
  NOR2_X1 prince_rounds_constant_MUX_U48 ( .A1(prince_rounds_constant_MUX_n13), 
        .A2(prince_rounds_constant_MUX_n26), .ZN(
        prince_rounds_constant_MUX_n38) );
  INV_X1 prince_rounds_constant_MUX_U47 ( .A(prince_rounds_constant_MUX_n24), 
        .ZN(prince_rounds_constant_MUX_n13) );
  NAND2_X1 prince_rounds_constant_MUX_U46 ( .A1(prince_rounds_constant_MUX_n18), .A2(prince_rounds_constant_MUX_n40), .ZN(prince_rounds_round_Constant[24])
         );
  AOI211_X1 prince_rounds_constant_MUX_U45 ( .C1(
        prince_rounds_constant_MUX_n20), .C2(prince_rounds_constant_MUX_n19), 
        .A(prince_rounds_constant_MUX_n12), .B(prince_rounds_constant_MUX_n11), 
        .ZN(prince_rounds_constant_MUX_n18) );
  INV_X1 prince_rounds_constant_MUX_U44 ( .A(prince_rounds_constant_MUX_n42), 
        .ZN(prince_rounds_constant_MUX_n11) );
  NAND2_X1 prince_rounds_constant_MUX_U43 ( .A1(prince_rounds_constant_MUX_n34), .A2(prince_rounds_constant_MUX_n32), .ZN(prince_rounds_round_Constant[22])
         );
  NAND2_X1 prince_rounds_constant_MUX_U42 ( .A1(prince_rounds_constant_MUX_n10), .A2(prince_rounds_constant_MUX_n20), .ZN(prince_rounds_constant_MUX_n32) );
  NOR2_X1 prince_rounds_constant_MUX_U41 ( .A1(prince_rounds_constant_MUX_n15), 
        .A2(prince_rounds_constant_MUX_n14), .ZN(
        prince_rounds_constant_MUX_n20) );
  AND2_X1 prince_rounds_constant_MUX_U40 ( .A1(prince_rounds_constant_MUX_n41), 
        .A2(prince_rounds_constant_MUX_n33), .ZN(
        prince_rounds_constant_MUX_n34) );
  NAND3_X1 prince_rounds_constant_MUX_U39 ( .A1(prince_rounds_constant_MUX_n33), .A2(prince_rounds_constant_MUX_n36), .A3(prince_rounds_constant_MUX_n40), 
        .ZN(prince_rounds_round_Constant[21]) );
  NAND3_X1 prince_rounds_constant_MUX_U38 ( .A1(prince_rounds_constant_MUX_n15), .A2(prince_rounds_constant_MUX_n16), .A3(prince_rounds_constant_MUX_n19), 
        .ZN(prince_rounds_constant_MUX_n40) );
  AND2_X1 prince_rounds_constant_MUX_U37 ( .A1(prince_rounds_constant_MUX_n42), 
        .A2(prince_rounds_constant_MUX_n21), .ZN(
        prince_rounds_constant_MUX_n33) );
  NAND2_X1 prince_rounds_constant_MUX_U36 ( .A1(prince_rounds_constant_MUX_n9), 
        .A2(prince_rounds_constant_MUX_n16), .ZN(
        prince_rounds_constant_MUX_n21) );
  AOI21_X1 prince_rounds_constant_MUX_U35 ( .B1(prince_rounds_constant_MUX_n10), .B2(prince_rounds_constant_MUX_n17), .A(prince_rounds_constant_MUX_n8), .ZN(
        prince_rounds_constant_MUX_n42) );
  NAND2_X1 prince_rounds_constant_MUX_U34 ( .A1(prince_rounds_constant_MUX_n36), .A2(prince_rounds_constant_MUX_n44), .ZN(prince_rounds_round_Constant[19])
         );
  AOI22_X1 prince_rounds_constant_MUX_U33 ( .A1(prince_rounds_constant_MUX_n10), .A2(prince_rounds_constant_MUX_n12), .B1(prince_rounds_constant_MUX_n7), 
        .B2(prince_rounds_constant_MUX_n9), .ZN(prince_rounds_constant_MUX_n36) );
  INV_X1 prince_rounds_constant_MUX_U32 ( .A(prince_rounds_constant_MUX_n6), 
        .ZN(prince_rounds_constant_MUX_n9) );
  NAND2_X1 prince_rounds_constant_MUX_U31 ( .A1(prince_rounds_constant_MUX_n41), .A2(prince_rounds_constant_MUX_n43), .ZN(prince_rounds_round_Constant[38])
         );
  NAND2_X1 prince_rounds_constant_MUX_U30 ( .A1(prince_rounds_constant_MUX_n15), .A2(prince_rounds_constant_MUX_n7), .ZN(prince_rounds_constant_MUX_n41) );
  INV_X1 prince_rounds_constant_MUX_U29 ( .A(prince_rounds_constant_MUX_n14), 
        .ZN(prince_rounds_constant_MUX_n7) );
  OAI21_X1 prince_rounds_constant_MUX_U28 ( .B1(prince_rounds_constant_MUX_n6), 
        .B2(prince_rounds_constant_MUX_n14), .A(prince_rounds_constant_MUX_n24), .ZN(prince_rounds_round_Constant[54]) );
  NAND2_X1 prince_rounds_constant_MUX_U27 ( .A1(prince_rounds_constant_MUX_n12), .A2(prince_rounds_constant_MUX_n19), .ZN(prince_rounds_constant_MUX_n24) );
  INV_X1 prince_rounds_constant_MUX_U26 ( .A(prince_rounds_constant_MUX_n45), 
        .ZN(prince_rounds_round_Constant[56]) );
  NOR2_X1 prince_rounds_constant_MUX_U25 ( .A1(
        prince_rounds_round_Constant[25]), .A2(prince_rounds_round_Constant[1]), .ZN(prince_rounds_constant_MUX_n45) );
  INV_X1 prince_rounds_constant_MUX_U24 ( .A(prince_rounds_constant_MUX_n23), 
        .ZN(prince_rounds_round_Constant[25]) );
  AOI21_X1 prince_rounds_constant_MUX_U23 ( .B1(prince_rounds_constant_MUX_n19), .B2(prince_rounds_constant_MUX_n17), .A(prince_rounds_constant_MUX_n8), .ZN(
        prince_rounds_constant_MUX_n23) );
  NOR3_X1 prince_rounds_constant_MUX_U22 ( .A1(prince_rounds_constant_MUX_n5), 
        .A2(prince_rounds_constant_MUX_n4), .A3(prince_rounds_constant_MUX_n6), 
        .ZN(prince_rounds_constant_MUX_n8) );
  NAND2_X1 prince_rounds_constant_MUX_U21 ( .A1(prince_rounds_constant_MUX_n10), .A2(prince_rounds_constant_MUX_n15), .ZN(prince_rounds_constant_MUX_n6) );
  INV_X1 prince_rounds_constant_MUX_U20 ( .A(prince_rounds_constant_MUX_n3), 
        .ZN(prince_rounds_constant_MUX_n5) );
  NOR2_X1 prince_rounds_constant_MUX_U19 ( .A1(prince_rounds_constant_MUX_n3), 
        .A2(prince_rounds_constant_MUX_n44), .ZN(
        prince_rounds_constant_MUX_n17) );
  NAND2_X1 prince_rounds_constant_MUX_U18 ( .A1(prince_rounds_constant_MUX_n4), 
        .A2(prince_rounds_constant_MUX_n2), .ZN(prince_rounds_constant_MUX_n44) );
  OAI21_X1 prince_rounds_constant_MUX_U17 ( .B1(prince_rounds_constant_MUX_n43), .B2(prince_rounds_constant_MUX_n19), .A(prince_rounds_constant_MUX_n1), .ZN(
        prince_rounds_round_Constant[1]) );
  INV_X1 prince_rounds_constant_MUX_U16 ( .A(prince_rounds_constant_MUX_n26), 
        .ZN(prince_rounds_constant_MUX_n1) );
  NOR3_X1 prince_rounds_constant_MUX_U15 ( .A1(prince_rounds_constant_MUX_n10), 
        .A2(prince_rounds_constant_MUX_n2), .A3(prince_rounds_constant_MUX_n14), .ZN(prince_rounds_constant_MUX_n26) );
  NAND2_X1 prince_rounds_constant_MUX_U14 ( .A1(prince_rounds_constant_MUX_n4), 
        .A2(prince_rounds_constant_MUX_n3), .ZN(prince_rounds_constant_MUX_n14) );
  INV_X1 prince_rounds_constant_MUX_U13 ( .A(prince_rounds_constant_MUX_n10), 
        .ZN(prince_rounds_constant_MUX_n19) );
  XOR2_X1 prince_rounds_constant_MUX_U12 ( .A(round_Signal[0]), .B(enc_dec), 
        .Z(prince_rounds_constant_MUX_n10) );
  INV_X1 prince_rounds_constant_MUX_U11 ( .A(prince_rounds_constant_MUX_n12), 
        .ZN(prince_rounds_constant_MUX_n43) );
  NOR2_X1 prince_rounds_constant_MUX_U10 ( .A1(prince_rounds_constant_MUX_n15), 
        .A2(prince_rounds_constant_MUX_n27), .ZN(
        prince_rounds_constant_MUX_n12) );
  INV_X1 prince_rounds_constant_MUX_U9 ( .A(prince_rounds_constant_MUX_n16), 
        .ZN(prince_rounds_constant_MUX_n27) );
  NOR2_X1 prince_rounds_constant_MUX_U8 ( .A1(prince_rounds_constant_MUX_n4), 
        .A2(prince_rounds_constant_MUX_n3), .ZN(prince_rounds_constant_MUX_n16) );
  XNOR2_X1 prince_rounds_constant_MUX_U7 ( .A(enc_dec), .B(round_Signal[3]), 
        .ZN(prince_rounds_constant_MUX_n3) );
  XOR2_X1 prince_rounds_constant_MUX_U6 ( .A(enc_dec), .B(round_Signal[2]), 
        .Z(prince_rounds_constant_MUX_n4) );
  XNOR2_X1 prince_rounds_constant_MUX_U5 ( .A(enc_dec), .B(round_Signal[1]), 
        .ZN(prince_rounds_constant_MUX_n2) );
  INV_X1 prince_rounds_constant_MUX_U4 ( .A(prince_rounds_constant_MUX_n2), 
        .ZN(prince_rounds_constant_MUX_n15) );
  AND2_X1 prince_rounds_constant_MUX_U3 ( .A1(prince_rounds_constant_MUX_n21), 
        .A2(prince_rounds_constant_MUX_n39), .ZN(
        prince_rounds_constant_MUX_n46) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_0_0_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_0_0_n3), .B(
        prince_rounds_round_Constant[53]), .ZN(
        prince_rounds_k1_XOR_round_Constant_0_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_0_0_U1 ( .A(1'b0), .B(Key1[0]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_0_0_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_0_1_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_0_1_n3), .B(
        prince_rounds_round_Constant[1]), .ZN(
        prince_rounds_k1_XOR_round_Constant_1_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_0_1_U1 ( .A(1'b0), .B(Key1[1]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_0_1_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_0_2_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_0_2_n3), .B(
        prince_rounds_round_Constant[34]), .ZN(
        prince_rounds_k1_XOR_round_Constant_2_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_0_2_U1 ( .A(1'b0), .B(Key1[2]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_0_2_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_0_3_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_0_3_n3), .B(
        prince_rounds_round_Constant[50]), .ZN(
        prince_rounds_k1_XOR_round_Constant_3_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_0_3_U1 ( .A(1'b0), .B(Key1[3]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_0_3_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_1_0_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_1_0_n3), .B(
        prince_rounds_round_Constant[4]), .ZN(
        prince_rounds_k1_XOR_round_Constant_4_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_1_0_U1 ( .A(1'b0), .B(Key1[4]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_1_0_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_1_1_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_1_1_n3), .B(
        prince_rounds_round_Constant[38]), .ZN(
        prince_rounds_k1_XOR_round_Constant_5_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_1_1_U1 ( .A(1'b0), .B(Key1[5]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_1_1_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_1_2_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_1_2_n3), .B(
        prince_rounds_round_Constant[33]), .ZN(
        prince_rounds_k1_XOR_round_Constant_6_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_1_2_U1 ( .A(1'b0), .B(Key1[6]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_1_2_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_1_3_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_1_3_n3), .B(
        prince_rounds_round_Constant[18]), .ZN(
        prince_rounds_k1_XOR_round_Constant_7_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_1_3_U1 ( .A(1'b0), .B(Key1[7]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_1_3_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_2_0_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_2_0_n3), .B(
        prince_rounds_round_Constant[8]), .ZN(
        prince_rounds_k1_XOR_round_Constant_8_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_2_0_U1 ( .A(1'b0), .B(Key1[8]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_2_0_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_2_1_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_2_1_n3), .B(
        prince_rounds_round_Constant[56]), .ZN(
        prince_rounds_k1_XOR_round_Constant_9_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_2_1_U1 ( .A(1'b0), .B(Key1[9]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_2_1_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_2_2_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_2_2_n3), .B(
        prince_rounds_round_Constant[59]), .ZN(
        prince_rounds_k1_XOR_round_Constant_10_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_2_2_U1 ( .A(1'b0), .B(Key1[10]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_2_2_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_2_3_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_2_3_n3), .B(
        prince_rounds_round_Constant[59]), .ZN(
        prince_rounds_k1_XOR_round_Constant_11_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_2_3_U1 ( .A(1'b0), .B(Key1[11]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_2_3_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_3_0_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_3_0_n3), .B(
        prince_rounds_round_Constant[37]), .ZN(
        prince_rounds_k1_XOR_round_Constant_12_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_3_0_U1 ( .A(1'b0), .B(Key1[12]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_3_0_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_3_1_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_3_1_n3), .B(
        prince_rounds_round_Constant[13]), .ZN(
        prince_rounds_k1_XOR_round_Constant_13_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_3_1_U1 ( .A(1'b0), .B(Key1[13]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_3_1_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_3_2_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_3_2_n3), .B(
        prince_rounds_round_Constant[14]), .ZN(
        prince_rounds_k1_XOR_round_Constant_14_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_3_2_U1 ( .A(1'b0), .B(Key1[14]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_3_2_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_3_3_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_3_3_n3), .B(1'b0), 
        .ZN(prince_rounds_k1_XOR_round_Constant_15_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_3_3_U1 ( .A(1'b0), .B(Key1[15]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_3_3_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_4_0_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_4_0_n3), .B(
        prince_rounds_round_Constant[61]), .ZN(
        prince_rounds_k1_XOR_round_Constant_16_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_4_0_U1 ( .A(1'b0), .B(Key1[16]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_4_0_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_4_1_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_4_1_n3), .B(
        prince_rounds_round_Constant[44]), .ZN(
        prince_rounds_k1_XOR_round_Constant_17_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_4_1_U1 ( .A(1'b0), .B(Key1[17]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_4_1_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_4_2_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_4_2_n3), .B(
        prince_rounds_round_Constant[18]), .ZN(
        prince_rounds_k1_XOR_round_Constant_18_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_4_2_U1 ( .A(1'b0), .B(Key1[18]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_4_2_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_4_3_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_4_3_n3), .B(
        prince_rounds_round_Constant[19]), .ZN(
        prince_rounds_k1_XOR_round_Constant_19_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_4_3_U1 ( .A(1'b0), .B(Key1[19]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_4_3_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_5_0_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_5_0_n3), .B(
        prince_rounds_round_Constant[37]), .ZN(
        prince_rounds_k1_XOR_round_Constant_20_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_5_0_U1 ( .A(1'b0), .B(Key1[20]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_5_0_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_5_1_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_5_1_n3), .B(
        prince_rounds_round_Constant[21]), .ZN(
        prince_rounds_k1_XOR_round_Constant_21_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_5_1_U1 ( .A(1'b0), .B(Key1[21]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_5_1_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_5_2_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_5_2_n3), .B(
        prince_rounds_round_Constant[22]), .ZN(
        prince_rounds_k1_XOR_round_Constant_22_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_5_2_U1 ( .A(1'b0), .B(Key1[22]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_5_2_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_5_3_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_5_3_n3), .B(
        prince_rounds_round_Constant[58]), .ZN(
        prince_rounds_k1_XOR_round_Constant_23_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_5_3_U1 ( .A(1'b0), .B(Key1[23]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_5_3_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_6_0_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_6_0_n3), .B(
        prince_rounds_round_Constant[24]), .ZN(
        prince_rounds_k1_XOR_round_Constant_24_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_6_0_U1 ( .A(1'b0), .B(Key1[24]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_6_0_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_6_1_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_6_1_n3), .B(
        prince_rounds_round_Constant[25]), .ZN(
        prince_rounds_k1_XOR_round_Constant_25_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_6_1_U1 ( .A(1'b0), .B(Key1[25]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_6_1_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_6_2_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_6_2_n3), .B(
        prince_rounds_round_Constant[59]), .ZN(
        prince_rounds_k1_XOR_round_Constant_26_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_6_2_U1 ( .A(1'b0), .B(Key1[26]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_6_2_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_6_3_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_6_3_n3), .B(
        prince_rounds_round_Constant[27]), .ZN(
        prince_rounds_k1_XOR_round_Constant_27_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_6_3_U1 ( .A(1'b0), .B(Key1[27]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_6_3_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_7_0_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_7_0_n3), .B(
        prince_rounds_round_Constant[38]), .ZN(
        prince_rounds_k1_XOR_round_Constant_28_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_7_0_U1 ( .A(1'b0), .B(Key1[28]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_7_0_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_7_1_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_7_1_n3), .B(
        prince_rounds_round_Constant[29]), .ZN(
        prince_rounds_k1_XOR_round_Constant_29_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_7_1_U1 ( .A(1'b0), .B(Key1[29]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_7_1_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_7_2_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_7_2_n3), .B(
        prince_rounds_round_Constant[36]), .ZN(
        prince_rounds_k1_XOR_round_Constant_30_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_7_2_U1 ( .A(1'b0), .B(Key1[30]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_7_2_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_7_3_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_7_3_n3), .B(
        prince_rounds_round_Constant[36]), .ZN(
        prince_rounds_k1_XOR_round_Constant_31_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_7_3_U1 ( .A(1'b0), .B(Key1[31]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_7_3_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_8_0_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_8_0_n3), .B(
        prince_rounds_round_Constant[32]), .ZN(
        prince_rounds_k1_XOR_round_Constant_32_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_8_0_U1 ( .A(1'b0), .B(Key1[32]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_8_0_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_8_1_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_8_1_n3), .B(
        prince_rounds_round_Constant[33]), .ZN(
        prince_rounds_k1_XOR_round_Constant_33_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_8_1_U1 ( .A(1'b0), .B(Key1[33]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_8_1_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_8_2_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_8_2_n3), .B(
        prince_rounds_round_Constant[34]), .ZN(
        prince_rounds_k1_XOR_round_Constant_34_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_8_2_U1 ( .A(1'b0), .B(Key1[34]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_8_2_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_8_3_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_8_3_n3), .B(
        prince_rounds_round_Constant[41]), .ZN(
        prince_rounds_k1_XOR_round_Constant_35_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_8_3_U1 ( .A(1'b0), .B(Key1[35]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_8_3_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_9_0_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_9_0_n3), .B(
        prince_rounds_round_Constant[36]), .ZN(
        prince_rounds_k1_XOR_round_Constant_36_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_9_0_U1 ( .A(1'b0), .B(Key1[36]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_9_0_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_9_1_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_9_1_n3), .B(
        prince_rounds_round_Constant[37]), .ZN(
        prince_rounds_k1_XOR_round_Constant_37_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_9_1_U1 ( .A(1'b0), .B(Key1[37]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_9_1_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_9_2_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_9_2_n3), .B(
        prince_rounds_round_Constant[38]), .ZN(
        prince_rounds_k1_XOR_round_Constant_38_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_9_2_U1 ( .A(1'b0), .B(Key1[38]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_9_2_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_9_3_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_9_3_n3), .B(
        prince_rounds_round_Constant[39]), .ZN(
        prince_rounds_k1_XOR_round_Constant_39_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_9_3_U1 ( .A(1'b0), .B(Key1[39]), .ZN(prince_rounds_k1_XOR_round_Constant_module_XORInst_9_3_n3)
         );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_10_0_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_10_0_n3), .B(
        prince_rounds_round_Constant[62]), .ZN(
        prince_rounds_k1_XOR_round_Constant_40_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_10_0_U1 ( .A(
        1'b0), .B(Key1[40]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_10_0_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_10_1_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_10_1_n3), .B(
        prince_rounds_round_Constant[41]), .ZN(
        prince_rounds_k1_XOR_round_Constant_41_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_10_1_U1 ( .A(
        1'b0), .B(Key1[41]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_10_1_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_10_2_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_10_2_n3), .B(
        prince_rounds_round_Constant[54]), .ZN(
        prince_rounds_k1_XOR_round_Constant_42_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_10_2_U1 ( .A(
        1'b0), .B(Key1[42]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_10_2_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_10_3_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_10_3_n3), .B(
        prince_rounds_round_Constant[43]), .ZN(
        prince_rounds_k1_XOR_round_Constant_43_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_10_3_U1 ( .A(
        1'b0), .B(Key1[43]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_10_3_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_11_0_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_11_0_n3), .B(
        prince_rounds_round_Constant[44]), .ZN(
        prince_rounds_k1_XOR_round_Constant_44_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_11_0_U1 ( .A(
        1'b0), .B(Key1[44]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_11_0_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_11_1_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_11_1_n3), .B(
        prince_rounds_round_Constant[45]), .ZN(
        prince_rounds_k1_XOR_round_Constant_45_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_11_1_U1 ( .A(
        1'b0), .B(Key1[45]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_11_1_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_11_2_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_11_2_n3), .B(
        prince_rounds_round_Constant[59]), .ZN(
        prince_rounds_k1_XOR_round_Constant_46_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_11_2_U1 ( .A(
        1'b0), .B(Key1[46]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_11_2_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_11_3_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_11_3_n3), .B(
        prince_rounds_round_Constant[47]), .ZN(
        prince_rounds_k1_XOR_round_Constant_47_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_11_3_U1 ( .A(
        1'b0), .B(Key1[47]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_11_3_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_12_0_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_12_0_n3), .B(
        prince_rounds_round_Constant[48]), .ZN(
        prince_rounds_k1_XOR_round_Constant_48_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_12_0_U1 ( .A(
        1'b0), .B(Key1[48]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_12_0_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_12_1_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_12_1_n3), .B(
        prince_rounds_round_Constant[49]), .ZN(
        prince_rounds_k1_XOR_round_Constant_49_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_12_1_U1 ( .A(
        1'b0), .B(Key1[49]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_12_1_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_12_2_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_12_2_n3), .B(
        prince_rounds_round_Constant[50]), .ZN(
        prince_rounds_k1_XOR_round_Constant_50_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_12_2_U1 ( .A(
        1'b0), .B(Key1[50]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_12_2_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_12_3_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_12_3_n3), .B(
        prince_rounds_round_Constant[51]), .ZN(
        prince_rounds_k1_XOR_round_Constant_51_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_12_3_U1 ( .A(
        1'b0), .B(Key1[51]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_12_3_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_13_0_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_13_0_n3), .B(
        prince_rounds_round_Constant[60]), .ZN(
        prince_rounds_k1_XOR_round_Constant_52_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_13_0_U1 ( .A(
        1'b0), .B(Key1[52]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_13_0_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_13_1_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_13_1_n3), .B(
        prince_rounds_round_Constant[53]), .ZN(
        prince_rounds_k1_XOR_round_Constant_53_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_13_1_U1 ( .A(
        1'b0), .B(Key1[53]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_13_1_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_13_2_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_13_2_n3), .B(
        prince_rounds_round_Constant[54]), .ZN(
        prince_rounds_k1_XOR_round_Constant_54_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_13_2_U1 ( .A(
        1'b0), .B(Key1[54]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_13_2_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_13_3_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_13_3_n3), .B(
        prince_rounds_round_Constant[55]), .ZN(
        prince_rounds_k1_XOR_round_Constant_55_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_13_3_U1 ( .A(
        1'b0), .B(Key1[55]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_13_3_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_14_0_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_14_0_n3), .B(
        prince_rounds_round_Constant[56]), .ZN(
        prince_rounds_k1_XOR_round_Constant_56_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_14_0_U1 ( .A(
        1'b0), .B(Key1[56]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_14_0_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_14_1_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_14_1_n3), .B(
        prince_rounds_round_Constant[60]), .ZN(
        prince_rounds_k1_XOR_round_Constant_57_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_14_1_U1 ( .A(
        1'b0), .B(Key1[57]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_14_1_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_14_2_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_14_2_n3), .B(
        prince_rounds_round_Constant[58]), .ZN(
        prince_rounds_k1_XOR_round_Constant_58_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_14_2_U1 ( .A(
        1'b0), .B(Key1[58]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_14_2_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_14_3_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_14_3_n3), .B(
        prince_rounds_round_Constant[59]), .ZN(
        prince_rounds_k1_XOR_round_Constant_59_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_14_3_U1 ( .A(
        1'b0), .B(Key1[59]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_14_3_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_15_0_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_15_0_n3), .B(
        prince_rounds_round_Constant[60]), .ZN(
        prince_rounds_k1_XOR_round_Constant_60_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_15_0_U1 ( .A(
        1'b0), .B(Key1[60]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_15_0_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_15_1_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_15_1_n3), .B(
        prince_rounds_round_Constant[61]), .ZN(
        prince_rounds_k1_XOR_round_Constant_61_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_15_1_U1 ( .A(
        1'b0), .B(Key1[61]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_15_1_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_15_2_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_15_2_n3), .B(
        prince_rounds_round_Constant[62]), .ZN(
        prince_rounds_k1_XOR_round_Constant_62_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_15_2_U1 ( .A(
        1'b0), .B(Key1[62]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_15_2_n3) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_15_3_U2 ( .A(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_15_3_n3), .B(
        prince_rounds_round_Constant[63]), .ZN(
        prince_rounds_k1_XOR_round_Constant_63_) );
  XNOR2_X1 prince_rounds_k1_XOR_round_Constant_module_XORInst_15_3_U1 ( .A(
        1'b0), .B(Key1[63]), .ZN(
        prince_rounds_k1_XOR_round_Constant_module_XORInst_15_3_n3) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_0_U1 ( .A(
        prince_rounds_mul_result_s1[0]), .B(prince_SR_Inv_Result_s1[0]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[48]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_1_U1 ( .A(
        prince_rounds_mul_result_s1[1]), .B(prince_SR_Inv_Result_s1[1]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[49]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_2_U1 ( .A(
        prince_rounds_mul_result_s1[2]), .B(prince_SR_Inv_Result_s1[2]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[50]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_3_U1 ( .A(
        prince_rounds_mul_result_s1[3]), .B(prince_SR_Inv_Result_s1[3]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[51]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_4_U1 ( .A(
        prince_rounds_mul_result_s1[4]), .B(prince_SR_Inv_Result_s1[4]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[36]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_5_U1 ( .A(
        prince_rounds_mul_result_s1[5]), .B(prince_SR_Inv_Result_s1[5]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[37]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_6_U1 ( .A(
        prince_rounds_mul_result_s1[6]), .B(prince_SR_Inv_Result_s1[6]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[38]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_7_U1 ( .A(
        prince_rounds_mul_result_s1[7]), .B(prince_SR_Inv_Result_s1[7]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[39]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_8_U1 ( .A(
        prince_rounds_mul_result_s1[8]), .B(prince_SR_Inv_Result_s1[8]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[24]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_9_U1 ( .A(
        prince_rounds_mul_result_s1[9]), .B(prince_SR_Inv_Result_s1[9]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[25]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_10_U1 ( .A(
        prince_rounds_mul_result_s1[10]), .B(prince_SR_Inv_Result_s1[10]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[26]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_11_U1 ( .A(
        prince_rounds_mul_result_s1[11]), .B(prince_SR_Inv_Result_s1[11]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[27]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_12_U1 ( .A(
        prince_rounds_mul_result_s1[12]), .B(prince_SR_Inv_Result_s1[12]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[12]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_13_U1 ( .A(
        prince_rounds_mul_result_s1[13]), .B(prince_SR_Inv_Result_s1[13]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[13]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_14_U1 ( .A(
        prince_rounds_mul_result_s1[14]), .B(prince_SR_Inv_Result_s1[14]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[14]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_15_U1 ( .A(
        prince_rounds_mul_result_s1[15]), .B(prince_SR_Inv_Result_s1[15]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[15]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_16_U1 ( .A(
        prince_rounds_mul_result_s1[16]), .B(prince_SR_Inv_Result_s1[16]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[0]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_17_U1 ( .A(
        prince_rounds_mul_result_s1[17]), .B(prince_SR_Inv_Result_s1[17]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[1]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_18_U1 ( .A(
        prince_rounds_mul_result_s1[18]), .B(prince_SR_Inv_Result_s1[18]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[2]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_19_U1 ( .A(
        prince_rounds_mul_result_s1[19]), .B(prince_SR_Inv_Result_s1[19]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[3]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_20_U1 ( .A(
        prince_rounds_mul_result_s1[20]), .B(prince_SR_Inv_Result_s1[20]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[52]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_21_U1 ( .A(
        prince_rounds_mul_result_s1[21]), .B(prince_SR_Inv_Result_s1[21]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[53]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_22_U1 ( .A(
        prince_rounds_mul_result_s1[22]), .B(prince_SR_Inv_Result_s1[22]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[54]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_23_U1 ( .A(
        prince_rounds_mul_result_s1[23]), .B(prince_SR_Inv_Result_s1[23]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[55]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_24_U1 ( .A(
        prince_rounds_mul_result_s1[24]), .B(prince_SR_Inv_Result_s1[24]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[40]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_25_U1 ( .A(
        prince_rounds_mul_result_s1[25]), .B(prince_SR_Inv_Result_s1[25]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[41]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_26_U1 ( .A(
        prince_rounds_mul_result_s1[26]), .B(prince_SR_Inv_Result_s1[26]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[42]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_27_U1 ( .A(
        prince_rounds_mul_result_s1[27]), .B(prince_SR_Inv_Result_s1[27]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[43]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_28_U1 ( .A(
        prince_rounds_mul_result_s1[28]), .B(prince_SR_Inv_Result_s1[28]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[28]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_29_U1 ( .A(
        prince_rounds_mul_result_s1[29]), .B(prince_SR_Inv_Result_s1[29]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[29]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_30_U1 ( .A(
        prince_rounds_mul_result_s1[30]), .B(prince_SR_Inv_Result_s1[30]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[30]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_31_U1 ( .A(
        prince_rounds_mul_result_s1[31]), .B(prince_SR_Inv_Result_s1[31]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[31]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_32_U1 ( .A(
        prince_rounds_mul_result_s1[32]), .B(prince_SR_Inv_Result_s1[32]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[16]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_33_U1 ( .A(
        prince_rounds_mul_result_s1[33]), .B(prince_SR_Inv_Result_s1[33]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[17]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_34_U1 ( .A(
        prince_rounds_mul_result_s1[34]), .B(prince_SR_Inv_Result_s1[34]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[18]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_35_U1 ( .A(
        prince_rounds_mul_result_s1[35]), .B(prince_SR_Inv_Result_s1[35]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[19]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_36_U1 ( .A(
        prince_rounds_mul_result_s1[36]), .B(prince_SR_Inv_Result_s1[36]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[4]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_37_U1 ( .A(
        prince_rounds_mul_result_s1[37]), .B(prince_SR_Inv_Result_s1[37]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[5]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_38_U1 ( .A(
        prince_rounds_mul_result_s1[38]), .B(prince_SR_Inv_Result_s1[38]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[6]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_39_U1 ( .A(
        prince_rounds_mul_result_s1[39]), .B(prince_SR_Inv_Result_s1[39]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[7]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_40_U1 ( .A(
        prince_rounds_mul_result_s1[40]), .B(prince_SR_Inv_Result_s1[40]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[56]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_41_U1 ( .A(
        prince_rounds_mul_result_s1[41]), .B(prince_SR_Inv_Result_s1[41]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[57]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_42_U1 ( .A(
        prince_rounds_mul_result_s1[42]), .B(prince_SR_Inv_Result_s1[42]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[58]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_43_U1 ( .A(
        prince_rounds_mul_result_s1[43]), .B(prince_SR_Inv_Result_s1[43]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[59]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_44_U1 ( .A(
        prince_rounds_mul_result_s1[44]), .B(prince_SR_Inv_Result_s1[44]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[44]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_45_U1 ( .A(
        prince_rounds_mul_result_s1[45]), .B(prince_SR_Inv_Result_s1[45]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[45]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_46_U1 ( .A(
        prince_rounds_mul_result_s1[46]), .B(prince_SR_Inv_Result_s1[46]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[46]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_47_U1 ( .A(
        prince_rounds_mul_result_s1[47]), .B(prince_SR_Inv_Result_s1[47]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[47]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_48_U1 ( .A(
        prince_rounds_mul_result_s1[48]), .B(prince_SR_Inv_Result_s1[48]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[32]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_49_U1 ( .A(
        prince_rounds_mul_result_s1[49]), .B(prince_SR_Inv_Result_s1[49]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[33]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_50_U1 ( .A(
        prince_rounds_mul_result_s1[50]), .B(prince_SR_Inv_Result_s1[50]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[34]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_51_U1 ( .A(
        prince_rounds_mul_result_s1[51]), .B(prince_SR_Inv_Result_s1[51]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[35]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_52_U1 ( .A(
        prince_rounds_mul_result_s1[52]), .B(prince_SR_Inv_Result_s1[52]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[20]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_53_U1 ( .A(
        prince_rounds_mul_result_s1[53]), .B(prince_SR_Inv_Result_s1[53]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[21]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_54_U1 ( .A(
        prince_rounds_mul_result_s1[54]), .B(prince_SR_Inv_Result_s1[54]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[22]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_55_U1 ( .A(
        prince_rounds_mul_result_s1[55]), .B(prince_SR_Inv_Result_s1[55]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[23]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_56_U1 ( .A(
        prince_rounds_mul_result_s1[56]), .B(prince_SR_Inv_Result_s1[56]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[8]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_57_U1 ( .A(
        prince_rounds_mul_result_s1[57]), .B(prince_SR_Inv_Result_s1[57]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[9]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_58_U1 ( .A(
        prince_rounds_mul_result_s1[58]), .B(prince_SR_Inv_Result_s1[58]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[10]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_59_U1 ( .A(
        prince_rounds_mul_result_s1[59]), .B(prince_SR_Inv_Result_s1[59]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[11]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_60_U1 ( .A(
        prince_rounds_mul_result_s1[60]), .B(prince_SR_Inv_Result_s1[60]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[60]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_61_U1 ( .A(
        prince_rounds_mul_result_s1[61]), .B(prince_SR_Inv_Result_s1[61]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[61]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_62_U1 ( .A(
        prince_rounds_mul_result_s1[62]), .B(prince_SR_Inv_Result_s1[62]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[62]) );
  MUX2_X1 prince_rounds_InputMUX1_MUXInst_63_U1 ( .A(
        prince_rounds_mul_result_s1[63]), .B(prince_SR_Inv_Result_s1[63]), .S(
        reset), .Z(prince_rounds_SR_Result_s1[63]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_0_U1 ( .A(
        prince_rounds_mul_result_s2[0]), .B(prince_SR_Inv_Result_s2[0]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[48]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_1_U1 ( .A(
        prince_rounds_mul_result_s2[1]), .B(prince_SR_Inv_Result_s2[1]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[49]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_2_U1 ( .A(
        prince_rounds_mul_result_s2[2]), .B(prince_SR_Inv_Result_s2[2]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[50]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_3_U1 ( .A(
        prince_rounds_mul_result_s2[3]), .B(prince_SR_Inv_Result_s2[3]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[51]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_4_U1 ( .A(
        prince_rounds_mul_result_s2[4]), .B(prince_SR_Inv_Result_s2[4]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[36]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_5_U1 ( .A(
        prince_rounds_mul_result_s2[5]), .B(prince_SR_Inv_Result_s2[5]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[37]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_6_U1 ( .A(
        prince_rounds_mul_result_s2[6]), .B(prince_SR_Inv_Result_s2[6]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[38]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_7_U1 ( .A(
        prince_rounds_mul_result_s2[7]), .B(prince_SR_Inv_Result_s2[7]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[39]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_8_U1 ( .A(
        prince_rounds_mul_result_s2[8]), .B(prince_SR_Inv_Result_s2[8]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[24]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_9_U1 ( .A(
        prince_rounds_mul_result_s2[9]), .B(prince_SR_Inv_Result_s2[9]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[25]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_10_U1 ( .A(
        prince_rounds_mul_result_s2[10]), .B(prince_SR_Inv_Result_s2[10]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[26]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_11_U1 ( .A(
        prince_rounds_mul_result_s2[11]), .B(prince_SR_Inv_Result_s2[11]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[27]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_12_U1 ( .A(
        prince_rounds_mul_result_s2[12]), .B(prince_SR_Inv_Result_s2[12]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[12]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_13_U1 ( .A(
        prince_rounds_mul_result_s2[13]), .B(prince_SR_Inv_Result_s2[13]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[13]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_14_U1 ( .A(
        prince_rounds_mul_result_s2[14]), .B(prince_SR_Inv_Result_s2[14]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[14]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_15_U1 ( .A(
        prince_rounds_mul_result_s2[15]), .B(prince_SR_Inv_Result_s2[15]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[15]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_16_U1 ( .A(
        prince_rounds_mul_result_s2[16]), .B(prince_SR_Inv_Result_s2[16]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[0]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_17_U1 ( .A(
        prince_rounds_mul_result_s2[17]), .B(prince_SR_Inv_Result_s2[17]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[1]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_18_U1 ( .A(
        prince_rounds_mul_result_s2[18]), .B(prince_SR_Inv_Result_s2[18]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[2]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_19_U1 ( .A(
        prince_rounds_mul_result_s2[19]), .B(prince_SR_Inv_Result_s2[19]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[3]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_20_U1 ( .A(
        prince_rounds_mul_result_s2[20]), .B(prince_SR_Inv_Result_s2[20]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[52]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_21_U1 ( .A(
        prince_rounds_mul_result_s2[21]), .B(prince_SR_Inv_Result_s2[21]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[53]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_22_U1 ( .A(
        prince_rounds_mul_result_s2[22]), .B(prince_SR_Inv_Result_s2[22]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[54]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_23_U1 ( .A(
        prince_rounds_mul_result_s2[23]), .B(prince_SR_Inv_Result_s2[23]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[55]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_24_U1 ( .A(
        prince_rounds_mul_result_s2[24]), .B(prince_SR_Inv_Result_s2[24]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[40]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_25_U1 ( .A(
        prince_rounds_mul_result_s2[25]), .B(prince_SR_Inv_Result_s2[25]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[41]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_26_U1 ( .A(
        prince_rounds_mul_result_s2[26]), .B(prince_SR_Inv_Result_s2[26]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[42]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_27_U1 ( .A(
        prince_rounds_mul_result_s2[27]), .B(prince_SR_Inv_Result_s2[27]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[43]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_28_U1 ( .A(
        prince_rounds_mul_result_s2[28]), .B(prince_SR_Inv_Result_s2[28]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[28]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_29_U1 ( .A(
        prince_rounds_mul_result_s2[29]), .B(prince_SR_Inv_Result_s2[29]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[29]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_30_U1 ( .A(
        prince_rounds_mul_result_s2[30]), .B(prince_SR_Inv_Result_s2[30]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[30]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_31_U1 ( .A(
        prince_rounds_mul_result_s2[31]), .B(prince_SR_Inv_Result_s2[31]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[31]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_32_U1 ( .A(
        prince_rounds_mul_result_s2[32]), .B(prince_SR_Inv_Result_s2[32]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[16]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_33_U1 ( .A(
        prince_rounds_mul_result_s2[33]), .B(prince_SR_Inv_Result_s2[33]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[17]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_34_U1 ( .A(
        prince_rounds_mul_result_s2[34]), .B(prince_SR_Inv_Result_s2[34]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[18]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_35_U1 ( .A(
        prince_rounds_mul_result_s2[35]), .B(prince_SR_Inv_Result_s2[35]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[19]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_36_U1 ( .A(
        prince_rounds_mul_result_s2[36]), .B(prince_SR_Inv_Result_s2[36]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[4]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_37_U1 ( .A(
        prince_rounds_mul_result_s2[37]), .B(prince_SR_Inv_Result_s2[37]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[5]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_38_U1 ( .A(
        prince_rounds_mul_result_s2[38]), .B(prince_SR_Inv_Result_s2[38]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[6]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_39_U1 ( .A(
        prince_rounds_mul_result_s2[39]), .B(prince_SR_Inv_Result_s2[39]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[7]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_40_U1 ( .A(
        prince_rounds_mul_result_s2[40]), .B(prince_SR_Inv_Result_s2[40]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[56]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_41_U1 ( .A(
        prince_rounds_mul_result_s2[41]), .B(prince_SR_Inv_Result_s2[41]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[57]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_42_U1 ( .A(
        prince_rounds_mul_result_s2[42]), .B(prince_SR_Inv_Result_s2[42]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[58]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_43_U1 ( .A(
        prince_rounds_mul_result_s2[43]), .B(prince_SR_Inv_Result_s2[43]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[59]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_44_U1 ( .A(
        prince_rounds_mul_result_s2[44]), .B(prince_SR_Inv_Result_s2[44]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[44]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_45_U1 ( .A(
        prince_rounds_mul_result_s2[45]), .B(prince_SR_Inv_Result_s2[45]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[45]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_46_U1 ( .A(
        prince_rounds_mul_result_s2[46]), .B(prince_SR_Inv_Result_s2[46]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[46]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_47_U1 ( .A(
        prince_rounds_mul_result_s2[47]), .B(prince_SR_Inv_Result_s2[47]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[47]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_48_U1 ( .A(
        prince_rounds_mul_result_s2[48]), .B(prince_SR_Inv_Result_s2[48]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[32]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_49_U1 ( .A(
        prince_rounds_mul_result_s2[49]), .B(prince_SR_Inv_Result_s2[49]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[33]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_50_U1 ( .A(
        prince_rounds_mul_result_s2[50]), .B(prince_SR_Inv_Result_s2[50]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[34]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_51_U1 ( .A(
        prince_rounds_mul_result_s2[51]), .B(prince_SR_Inv_Result_s2[51]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[35]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_52_U1 ( .A(
        prince_rounds_mul_result_s2[52]), .B(prince_SR_Inv_Result_s2[52]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[20]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_53_U1 ( .A(
        prince_rounds_mul_result_s2[53]), .B(prince_SR_Inv_Result_s2[53]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[21]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_54_U1 ( .A(
        prince_rounds_mul_result_s2[54]), .B(prince_SR_Inv_Result_s2[54]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[22]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_55_U1 ( .A(
        prince_rounds_mul_result_s2[55]), .B(prince_SR_Inv_Result_s2[55]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[23]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_56_U1 ( .A(
        prince_rounds_mul_result_s2[56]), .B(prince_SR_Inv_Result_s2[56]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[8]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_57_U1 ( .A(
        prince_rounds_mul_result_s2[57]), .B(prince_SR_Inv_Result_s2[57]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[9]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_58_U1 ( .A(
        prince_rounds_mul_result_s2[58]), .B(prince_SR_Inv_Result_s2[58]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[10]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_59_U1 ( .A(
        prince_rounds_mul_result_s2[59]), .B(prince_SR_Inv_Result_s2[59]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[11]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_60_U1 ( .A(
        prince_rounds_mul_result_s2[60]), .B(prince_SR_Inv_Result_s2[60]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[60]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_61_U1 ( .A(
        prince_rounds_mul_result_s2[61]), .B(prince_SR_Inv_Result_s2[61]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[61]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_62_U1 ( .A(
        prince_rounds_mul_result_s2[62]), .B(prince_SR_Inv_Result_s2[62]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[62]) );
  MUX2_X1 prince_rounds_InputMUX2_MUXInst_63_U1 ( .A(
        prince_rounds_mul_result_s2[63]), .B(prince_SR_Inv_Result_s2[63]), .S(
        reset), .Z(prince_rounds_SR_Result_s2[63]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_0_U1 ( .A(
        prince_rounds_mul_result_s3[0]), .B(prince_SR_Inv_Result_s3[0]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[48]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_1_U1 ( .A(
        prince_rounds_mul_result_s3[1]), .B(prince_SR_Inv_Result_s3[1]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[49]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_2_U1 ( .A(
        prince_rounds_mul_result_s3[2]), .B(prince_SR_Inv_Result_s3[2]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[50]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_3_U1 ( .A(
        prince_rounds_mul_result_s3[3]), .B(prince_SR_Inv_Result_s3[3]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[51]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_4_U1 ( .A(
        prince_rounds_mul_result_s3[4]), .B(prince_SR_Inv_Result_s3[4]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[36]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_5_U1 ( .A(
        prince_rounds_mul_result_s3[5]), .B(prince_SR_Inv_Result_s3[5]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[37]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_6_U1 ( .A(
        prince_rounds_mul_result_s3[6]), .B(prince_SR_Inv_Result_s3[6]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[38]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_7_U1 ( .A(
        prince_rounds_mul_result_s3[7]), .B(prince_SR_Inv_Result_s3[7]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[39]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_8_U1 ( .A(
        prince_rounds_mul_result_s3[8]), .B(prince_SR_Inv_Result_s3[8]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[24]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_9_U1 ( .A(
        prince_rounds_mul_result_s3[9]), .B(prince_SR_Inv_Result_s3[9]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[25]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_10_U1 ( .A(
        prince_rounds_mul_result_s3[10]), .B(prince_SR_Inv_Result_s3[10]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[26]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_11_U1 ( .A(
        prince_rounds_mul_result_s3[11]), .B(prince_SR_Inv_Result_s3[11]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[27]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_12_U1 ( .A(
        prince_rounds_mul_result_s3[12]), .B(prince_SR_Inv_Result_s3[12]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[12]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_13_U1 ( .A(
        prince_rounds_mul_result_s3[13]), .B(prince_SR_Inv_Result_s3[13]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[13]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_14_U1 ( .A(
        prince_rounds_mul_result_s3[14]), .B(prince_SR_Inv_Result_s3[14]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[14]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_15_U1 ( .A(
        prince_rounds_mul_result_s3[15]), .B(prince_SR_Inv_Result_s3[15]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[15]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_16_U1 ( .A(
        prince_rounds_mul_result_s3[16]), .B(prince_SR_Inv_Result_s3[16]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[0]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_17_U1 ( .A(
        prince_rounds_mul_result_s3[17]), .B(prince_SR_Inv_Result_s3[17]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[1]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_18_U1 ( .A(
        prince_rounds_mul_result_s3[18]), .B(prince_SR_Inv_Result_s3[18]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[2]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_19_U1 ( .A(
        prince_rounds_mul_result_s3[19]), .B(prince_SR_Inv_Result_s3[19]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[3]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_20_U1 ( .A(
        prince_rounds_mul_result_s3[20]), .B(prince_SR_Inv_Result_s3[20]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[52]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_21_U1 ( .A(
        prince_rounds_mul_result_s3[21]), .B(prince_SR_Inv_Result_s3[21]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[53]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_22_U1 ( .A(
        prince_rounds_mul_result_s3[22]), .B(prince_SR_Inv_Result_s3[22]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[54]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_23_U1 ( .A(
        prince_rounds_mul_result_s3[23]), .B(prince_SR_Inv_Result_s3[23]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[55]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_24_U1 ( .A(
        prince_rounds_mul_result_s3[24]), .B(prince_SR_Inv_Result_s3[24]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[40]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_25_U1 ( .A(
        prince_rounds_mul_result_s3[25]), .B(prince_SR_Inv_Result_s3[25]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[41]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_26_U1 ( .A(
        prince_rounds_mul_result_s3[26]), .B(prince_SR_Inv_Result_s3[26]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[42]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_27_U1 ( .A(
        prince_rounds_mul_result_s3[27]), .B(prince_SR_Inv_Result_s3[27]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[43]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_28_U1 ( .A(
        prince_rounds_mul_result_s3[28]), .B(prince_SR_Inv_Result_s3[28]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[28]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_29_U1 ( .A(
        prince_rounds_mul_result_s3[29]), .B(prince_SR_Inv_Result_s3[29]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[29]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_30_U1 ( .A(
        prince_rounds_mul_result_s3[30]), .B(prince_SR_Inv_Result_s3[30]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[30]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_31_U1 ( .A(
        prince_rounds_mul_result_s3[31]), .B(prince_SR_Inv_Result_s3[31]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[31]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_32_U1 ( .A(
        prince_rounds_mul_result_s3[32]), .B(prince_SR_Inv_Result_s3[32]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[16]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_33_U1 ( .A(
        prince_rounds_mul_result_s3[33]), .B(prince_SR_Inv_Result_s3[33]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[17]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_34_U1 ( .A(
        prince_rounds_mul_result_s3[34]), .B(prince_SR_Inv_Result_s3[34]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[18]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_35_U1 ( .A(
        prince_rounds_mul_result_s3[35]), .B(prince_SR_Inv_Result_s3[35]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[19]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_36_U1 ( .A(
        prince_rounds_mul_result_s3[36]), .B(prince_SR_Inv_Result_s3[36]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[4]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_37_U1 ( .A(
        prince_rounds_mul_result_s3[37]), .B(prince_SR_Inv_Result_s3[37]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[5]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_38_U1 ( .A(
        prince_rounds_mul_result_s3[38]), .B(prince_SR_Inv_Result_s3[38]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[6]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_39_U1 ( .A(
        prince_rounds_mul_result_s3[39]), .B(prince_SR_Inv_Result_s3[39]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[7]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_40_U1 ( .A(
        prince_rounds_mul_result_s3[40]), .B(prince_SR_Inv_Result_s3[40]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[56]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_41_U1 ( .A(
        prince_rounds_mul_result_s3[41]), .B(prince_SR_Inv_Result_s3[41]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[57]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_42_U1 ( .A(
        prince_rounds_mul_result_s3[42]), .B(prince_SR_Inv_Result_s3[42]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[58]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_43_U1 ( .A(
        prince_rounds_mul_result_s3[43]), .B(prince_SR_Inv_Result_s3[43]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[59]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_44_U1 ( .A(
        prince_rounds_mul_result_s3[44]), .B(prince_SR_Inv_Result_s3[44]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[44]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_45_U1 ( .A(
        prince_rounds_mul_result_s3[45]), .B(prince_SR_Inv_Result_s3[45]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[45]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_46_U1 ( .A(
        prince_rounds_mul_result_s3[46]), .B(prince_SR_Inv_Result_s3[46]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[46]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_47_U1 ( .A(
        prince_rounds_mul_result_s3[47]), .B(prince_SR_Inv_Result_s3[47]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[47]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_48_U1 ( .A(
        prince_rounds_mul_result_s3[48]), .B(prince_SR_Inv_Result_s3[48]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[32]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_49_U1 ( .A(
        prince_rounds_mul_result_s3[49]), .B(prince_SR_Inv_Result_s3[49]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[33]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_50_U1 ( .A(
        prince_rounds_mul_result_s3[50]), .B(prince_SR_Inv_Result_s3[50]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[34]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_51_U1 ( .A(
        prince_rounds_mul_result_s3[51]), .B(prince_SR_Inv_Result_s3[51]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[35]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_52_U1 ( .A(
        prince_rounds_mul_result_s3[52]), .B(prince_SR_Inv_Result_s3[52]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[20]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_53_U1 ( .A(
        prince_rounds_mul_result_s3[53]), .B(prince_SR_Inv_Result_s3[53]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[21]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_54_U1 ( .A(
        prince_rounds_mul_result_s3[54]), .B(prince_SR_Inv_Result_s3[54]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[22]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_55_U1 ( .A(
        prince_rounds_mul_result_s3[55]), .B(prince_SR_Inv_Result_s3[55]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[23]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_56_U1 ( .A(
        prince_rounds_mul_result_s3[56]), .B(prince_SR_Inv_Result_s3[56]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[8]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_57_U1 ( .A(
        prince_rounds_mul_result_s3[57]), .B(prince_SR_Inv_Result_s3[57]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[9]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_58_U1 ( .A(
        prince_rounds_mul_result_s3[58]), .B(prince_SR_Inv_Result_s3[58]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[10]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_59_U1 ( .A(
        prince_rounds_mul_result_s3[59]), .B(prince_SR_Inv_Result_s3[59]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[11]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_60_U1 ( .A(
        prince_rounds_mul_result_s3[60]), .B(prince_SR_Inv_Result_s3[60]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[60]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_61_U1 ( .A(
        prince_rounds_mul_result_s3[61]), .B(prince_SR_Inv_Result_s3[61]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[61]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_62_U1 ( .A(
        prince_rounds_mul_result_s3[62]), .B(prince_SR_Inv_Result_s3[62]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[62]) );
  MUX2_X1 prince_rounds_InputMUX3_MUXInst_63_U1 ( .A(
        prince_rounds_mul_result_s3[63]), .B(prince_SR_Inv_Result_s3[63]), .S(
        reset), .Z(prince_rounds_SR_Result_s3[63]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_0_0_U2 ( .A(
        prince_rounds_AddKey1_XORInst_0_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_0_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[0]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_0_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[0]), .ZN(
        prince_rounds_AddKey1_XORInst_0_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_0_1_U2 ( .A(
        prince_rounds_AddKey1_XORInst_0_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_1_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[1]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_0_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[1]), .ZN(
        prince_rounds_AddKey1_XORInst_0_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_0_2_U2 ( .A(
        prince_rounds_AddKey1_XORInst_0_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_2_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[2]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_0_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[2]), .ZN(
        prince_rounds_AddKey1_XORInst_0_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_0_3_U2 ( .A(
        prince_rounds_AddKey1_XORInst_0_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_3_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[3]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_0_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[3]), .ZN(
        prince_rounds_AddKey1_XORInst_0_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_1_0_U2 ( .A(
        prince_rounds_AddKey1_XORInst_1_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_4_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[4]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_1_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[4]), .ZN(
        prince_rounds_AddKey1_XORInst_1_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_1_1_U2 ( .A(
        prince_rounds_AddKey1_XORInst_1_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_5_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[5]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_1_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[5]), .ZN(
        prince_rounds_AddKey1_XORInst_1_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_1_2_U2 ( .A(
        prince_rounds_AddKey1_XORInst_1_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_6_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[6]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_1_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[6]), .ZN(
        prince_rounds_AddKey1_XORInst_1_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_1_3_U2 ( .A(
        prince_rounds_AddKey1_XORInst_1_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_7_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[7]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_1_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[7]), .ZN(
        prince_rounds_AddKey1_XORInst_1_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_2_0_U2 ( .A(
        prince_rounds_AddKey1_XORInst_2_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_8_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[8]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_2_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[8]), .ZN(
        prince_rounds_AddKey1_XORInst_2_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_2_1_U2 ( .A(
        prince_rounds_AddKey1_XORInst_2_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_9_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[9]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_2_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[9]), .ZN(
        prince_rounds_AddKey1_XORInst_2_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_2_2_U2 ( .A(
        prince_rounds_AddKey1_XORInst_2_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_10_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[10]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_2_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[10]), .ZN(
        prince_rounds_AddKey1_XORInst_2_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_2_3_U2 ( .A(
        prince_rounds_AddKey1_XORInst_2_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_11_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[11]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_2_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[11]), .ZN(
        prince_rounds_AddKey1_XORInst_2_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_3_0_U2 ( .A(
        prince_rounds_AddKey1_XORInst_3_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_12_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[12]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_3_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[12]), .ZN(
        prince_rounds_AddKey1_XORInst_3_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_3_1_U2 ( .A(
        prince_rounds_AddKey1_XORInst_3_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_13_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[13]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_3_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[13]), .ZN(
        prince_rounds_AddKey1_XORInst_3_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_3_2_U2 ( .A(
        prince_rounds_AddKey1_XORInst_3_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_14_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[14]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_3_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[14]), .ZN(
        prince_rounds_AddKey1_XORInst_3_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_3_3_U2 ( .A(
        prince_rounds_AddKey1_XORInst_3_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_15_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[15]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_3_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[15]), .ZN(
        prince_rounds_AddKey1_XORInst_3_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_4_0_U2 ( .A(
        prince_rounds_AddKey1_XORInst_4_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_16_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[16]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_4_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[16]), .ZN(
        prince_rounds_AddKey1_XORInst_4_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_4_1_U2 ( .A(
        prince_rounds_AddKey1_XORInst_4_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_17_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[17]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_4_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[17]), .ZN(
        prince_rounds_AddKey1_XORInst_4_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_4_2_U2 ( .A(
        prince_rounds_AddKey1_XORInst_4_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_18_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[18]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_4_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[18]), .ZN(
        prince_rounds_AddKey1_XORInst_4_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_4_3_U2 ( .A(
        prince_rounds_AddKey1_XORInst_4_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_19_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[19]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_4_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[19]), .ZN(
        prince_rounds_AddKey1_XORInst_4_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_5_0_U2 ( .A(
        prince_rounds_AddKey1_XORInst_5_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_20_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[20]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_5_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[20]), .ZN(
        prince_rounds_AddKey1_XORInst_5_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_5_1_U2 ( .A(
        prince_rounds_AddKey1_XORInst_5_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_21_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[21]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_5_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[21]), .ZN(
        prince_rounds_AddKey1_XORInst_5_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_5_2_U2 ( .A(
        prince_rounds_AddKey1_XORInst_5_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_22_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[22]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_5_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[22]), .ZN(
        prince_rounds_AddKey1_XORInst_5_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_5_3_U2 ( .A(
        prince_rounds_AddKey1_XORInst_5_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_23_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[23]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_5_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[23]), .ZN(
        prince_rounds_AddKey1_XORInst_5_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_6_0_U2 ( .A(
        prince_rounds_AddKey1_XORInst_6_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_24_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[24]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_6_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[24]), .ZN(
        prince_rounds_AddKey1_XORInst_6_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_6_1_U2 ( .A(
        prince_rounds_AddKey1_XORInst_6_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_25_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[25]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_6_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[25]), .ZN(
        prince_rounds_AddKey1_XORInst_6_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_6_2_U2 ( .A(
        prince_rounds_AddKey1_XORInst_6_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_26_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[26]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_6_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[26]), .ZN(
        prince_rounds_AddKey1_XORInst_6_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_6_3_U2 ( .A(
        prince_rounds_AddKey1_XORInst_6_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_27_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[27]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_6_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[27]), .ZN(
        prince_rounds_AddKey1_XORInst_6_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_7_0_U2 ( .A(
        prince_rounds_AddKey1_XORInst_7_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_28_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[28]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_7_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[28]), .ZN(
        prince_rounds_AddKey1_XORInst_7_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_7_1_U2 ( .A(
        prince_rounds_AddKey1_XORInst_7_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_29_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[29]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_7_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[29]), .ZN(
        prince_rounds_AddKey1_XORInst_7_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_7_2_U2 ( .A(
        prince_rounds_AddKey1_XORInst_7_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_30_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[30]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_7_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[30]), .ZN(
        prince_rounds_AddKey1_XORInst_7_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_7_3_U2 ( .A(
        prince_rounds_AddKey1_XORInst_7_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_31_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[31]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_7_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[31]), .ZN(
        prince_rounds_AddKey1_XORInst_7_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_8_0_U2 ( .A(
        prince_rounds_AddKey1_XORInst_8_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_32_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[32]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_8_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[32]), .ZN(
        prince_rounds_AddKey1_XORInst_8_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_8_1_U2 ( .A(
        prince_rounds_AddKey1_XORInst_8_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_33_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[33]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_8_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[33]), .ZN(
        prince_rounds_AddKey1_XORInst_8_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_8_2_U2 ( .A(
        prince_rounds_AddKey1_XORInst_8_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_34_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[34]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_8_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[34]), .ZN(
        prince_rounds_AddKey1_XORInst_8_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_8_3_U2 ( .A(
        prince_rounds_AddKey1_XORInst_8_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_35_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[35]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_8_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[35]), .ZN(
        prince_rounds_AddKey1_XORInst_8_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_9_0_U2 ( .A(
        prince_rounds_AddKey1_XORInst_9_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_36_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[36]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_9_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[36]), .ZN(
        prince_rounds_AddKey1_XORInst_9_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_9_1_U2 ( .A(
        prince_rounds_AddKey1_XORInst_9_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_37_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[37]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_9_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[37]), .ZN(
        prince_rounds_AddKey1_XORInst_9_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_9_2_U2 ( .A(
        prince_rounds_AddKey1_XORInst_9_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_38_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[38]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_9_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[38]), .ZN(
        prince_rounds_AddKey1_XORInst_9_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_9_3_U2 ( .A(
        prince_rounds_AddKey1_XORInst_9_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_39_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[39]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_9_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[39]), .ZN(
        prince_rounds_AddKey1_XORInst_9_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_10_0_U2 ( .A(
        prince_rounds_AddKey1_XORInst_10_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_40_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[40]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_10_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[40]), .ZN(
        prince_rounds_AddKey1_XORInst_10_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_10_1_U2 ( .A(
        prince_rounds_AddKey1_XORInst_10_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_41_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[41]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_10_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[41]), .ZN(
        prince_rounds_AddKey1_XORInst_10_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_10_2_U2 ( .A(
        prince_rounds_AddKey1_XORInst_10_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_42_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[42]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_10_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[42]), .ZN(
        prince_rounds_AddKey1_XORInst_10_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_10_3_U2 ( .A(
        prince_rounds_AddKey1_XORInst_10_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_43_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[43]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_10_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[43]), .ZN(
        prince_rounds_AddKey1_XORInst_10_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_11_0_U2 ( .A(
        prince_rounds_AddKey1_XORInst_11_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_44_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[44]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_11_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[44]), .ZN(
        prince_rounds_AddKey1_XORInst_11_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_11_1_U2 ( .A(
        prince_rounds_AddKey1_XORInst_11_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_45_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[45]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_11_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[45]), .ZN(
        prince_rounds_AddKey1_XORInst_11_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_11_2_U2 ( .A(
        prince_rounds_AddKey1_XORInst_11_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_46_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[46]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_11_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[46]), .ZN(
        prince_rounds_AddKey1_XORInst_11_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_11_3_U2 ( .A(
        prince_rounds_AddKey1_XORInst_11_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_47_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[47]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_11_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[47]), .ZN(
        prince_rounds_AddKey1_XORInst_11_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_12_0_U2 ( .A(
        prince_rounds_AddKey1_XORInst_12_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_48_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[48]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_12_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[48]), .ZN(
        prince_rounds_AddKey1_XORInst_12_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_12_1_U2 ( .A(
        prince_rounds_AddKey1_XORInst_12_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_49_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[49]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_12_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[49]), .ZN(
        prince_rounds_AddKey1_XORInst_12_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_12_2_U2 ( .A(
        prince_rounds_AddKey1_XORInst_12_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_50_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[50]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_12_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[50]), .ZN(
        prince_rounds_AddKey1_XORInst_12_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_12_3_U2 ( .A(
        prince_rounds_AddKey1_XORInst_12_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_51_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[51]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_12_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[51]), .ZN(
        prince_rounds_AddKey1_XORInst_12_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_13_0_U2 ( .A(
        prince_rounds_AddKey1_XORInst_13_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_52_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[52]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_13_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[52]), .ZN(
        prince_rounds_AddKey1_XORInst_13_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_13_1_U2 ( .A(
        prince_rounds_AddKey1_XORInst_13_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_53_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[53]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_13_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[53]), .ZN(
        prince_rounds_AddKey1_XORInst_13_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_13_2_U2 ( .A(
        prince_rounds_AddKey1_XORInst_13_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_54_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[54]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_13_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[54]), .ZN(
        prince_rounds_AddKey1_XORInst_13_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_13_3_U2 ( .A(
        prince_rounds_AddKey1_XORInst_13_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_55_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[55]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_13_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[55]), .ZN(
        prince_rounds_AddKey1_XORInst_13_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_14_0_U2 ( .A(
        prince_rounds_AddKey1_XORInst_14_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_56_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[56]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_14_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[56]), .ZN(
        prince_rounds_AddKey1_XORInst_14_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_14_1_U2 ( .A(
        prince_rounds_AddKey1_XORInst_14_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_57_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[57]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_14_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[57]), .ZN(
        prince_rounds_AddKey1_XORInst_14_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_14_2_U2 ( .A(
        prince_rounds_AddKey1_XORInst_14_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_58_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[58]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_14_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[58]), .ZN(
        prince_rounds_AddKey1_XORInst_14_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_14_3_U2 ( .A(
        prince_rounds_AddKey1_XORInst_14_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_59_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[59]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_14_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[59]), .ZN(
        prince_rounds_AddKey1_XORInst_14_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_15_0_U2 ( .A(
        prince_rounds_AddKey1_XORInst_15_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_60_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[60]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_15_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[60]), .ZN(
        prince_rounds_AddKey1_XORInst_15_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_15_1_U2 ( .A(
        prince_rounds_AddKey1_XORInst_15_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_61_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[61]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_15_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[61]), .ZN(
        prince_rounds_AddKey1_XORInst_15_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_15_2_U2 ( .A(
        prince_rounds_AddKey1_XORInst_15_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_62_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[62]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_15_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[62]), .ZN(
        prince_rounds_AddKey1_XORInst_15_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_15_3_U2 ( .A(
        prince_rounds_AddKey1_XORInst_15_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_63_), .ZN(
        prince_rounds_round_inputXORkeyRCON_s1[63]) );
  XNOR2_X1 prince_rounds_AddKey1_XORInst_15_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s1[63]), .ZN(
        prince_rounds_AddKey1_XORInst_15_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_0_0_U2 ( .A(
        prince_rounds_AddKey2_XORInst_0_0_n3), .B(Key2[0]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[0]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_0_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[0]), .ZN(
        prince_rounds_AddKey2_XORInst_0_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_0_1_U2 ( .A(
        prince_rounds_AddKey2_XORInst_0_1_n3), .B(Key2[1]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[1]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_0_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[1]), .ZN(
        prince_rounds_AddKey2_XORInst_0_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_0_2_U2 ( .A(
        prince_rounds_AddKey2_XORInst_0_2_n3), .B(Key2[2]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[2]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_0_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[2]), .ZN(
        prince_rounds_AddKey2_XORInst_0_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_0_3_U2 ( .A(
        prince_rounds_AddKey2_XORInst_0_3_n3), .B(Key2[3]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[3]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_0_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[3]), .ZN(
        prince_rounds_AddKey2_XORInst_0_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_1_0_U2 ( .A(
        prince_rounds_AddKey2_XORInst_1_0_n3), .B(Key2[4]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[4]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_1_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[4]), .ZN(
        prince_rounds_AddKey2_XORInst_1_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_1_1_U2 ( .A(
        prince_rounds_AddKey2_XORInst_1_1_n3), .B(Key2[5]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[5]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_1_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[5]), .ZN(
        prince_rounds_AddKey2_XORInst_1_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_1_2_U2 ( .A(
        prince_rounds_AddKey2_XORInst_1_2_n3), .B(Key2[6]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[6]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_1_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[6]), .ZN(
        prince_rounds_AddKey2_XORInst_1_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_1_3_U2 ( .A(
        prince_rounds_AddKey2_XORInst_1_3_n3), .B(Key2[7]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[7]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_1_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[7]), .ZN(
        prince_rounds_AddKey2_XORInst_1_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_2_0_U2 ( .A(
        prince_rounds_AddKey2_XORInst_2_0_n3), .B(Key2[8]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[8]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_2_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[8]), .ZN(
        prince_rounds_AddKey2_XORInst_2_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_2_1_U2 ( .A(
        prince_rounds_AddKey2_XORInst_2_1_n3), .B(Key2[9]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[9]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_2_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[9]), .ZN(
        prince_rounds_AddKey2_XORInst_2_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_2_2_U2 ( .A(
        prince_rounds_AddKey2_XORInst_2_2_n3), .B(Key2[10]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[10]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_2_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[10]), .ZN(
        prince_rounds_AddKey2_XORInst_2_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_2_3_U2 ( .A(
        prince_rounds_AddKey2_XORInst_2_3_n3), .B(Key2[11]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[11]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_2_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[11]), .ZN(
        prince_rounds_AddKey2_XORInst_2_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_3_0_U2 ( .A(
        prince_rounds_AddKey2_XORInst_3_0_n3), .B(Key2[12]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[12]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_3_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[12]), .ZN(
        prince_rounds_AddKey2_XORInst_3_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_3_1_U2 ( .A(
        prince_rounds_AddKey2_XORInst_3_1_n3), .B(Key2[13]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[13]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_3_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[13]), .ZN(
        prince_rounds_AddKey2_XORInst_3_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_3_2_U2 ( .A(
        prince_rounds_AddKey2_XORInst_3_2_n3), .B(Key2[14]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[14]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_3_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[14]), .ZN(
        prince_rounds_AddKey2_XORInst_3_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_3_3_U2 ( .A(
        prince_rounds_AddKey2_XORInst_3_3_n3), .B(Key2[15]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[15]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_3_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[15]), .ZN(
        prince_rounds_AddKey2_XORInst_3_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_4_0_U2 ( .A(
        prince_rounds_AddKey2_XORInst_4_0_n3), .B(Key2[16]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[16]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_4_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[16]), .ZN(
        prince_rounds_AddKey2_XORInst_4_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_4_1_U2 ( .A(
        prince_rounds_AddKey2_XORInst_4_1_n3), .B(Key2[17]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[17]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_4_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[17]), .ZN(
        prince_rounds_AddKey2_XORInst_4_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_4_2_U2 ( .A(
        prince_rounds_AddKey2_XORInst_4_2_n3), .B(Key2[18]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[18]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_4_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[18]), .ZN(
        prince_rounds_AddKey2_XORInst_4_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_4_3_U2 ( .A(
        prince_rounds_AddKey2_XORInst_4_3_n3), .B(Key2[19]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[19]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_4_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[19]), .ZN(
        prince_rounds_AddKey2_XORInst_4_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_5_0_U2 ( .A(
        prince_rounds_AddKey2_XORInst_5_0_n3), .B(Key2[20]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[20]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_5_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[20]), .ZN(
        prince_rounds_AddKey2_XORInst_5_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_5_1_U2 ( .A(
        prince_rounds_AddKey2_XORInst_5_1_n3), .B(Key2[21]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[21]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_5_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[21]), .ZN(
        prince_rounds_AddKey2_XORInst_5_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_5_2_U2 ( .A(
        prince_rounds_AddKey2_XORInst_5_2_n3), .B(Key2[22]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[22]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_5_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[22]), .ZN(
        prince_rounds_AddKey2_XORInst_5_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_5_3_U2 ( .A(
        prince_rounds_AddKey2_XORInst_5_3_n3), .B(Key2[23]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[23]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_5_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[23]), .ZN(
        prince_rounds_AddKey2_XORInst_5_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_6_0_U2 ( .A(
        prince_rounds_AddKey2_XORInst_6_0_n3), .B(Key2[24]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[24]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_6_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[24]), .ZN(
        prince_rounds_AddKey2_XORInst_6_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_6_1_U2 ( .A(
        prince_rounds_AddKey2_XORInst_6_1_n3), .B(Key2[25]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[25]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_6_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[25]), .ZN(
        prince_rounds_AddKey2_XORInst_6_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_6_2_U2 ( .A(
        prince_rounds_AddKey2_XORInst_6_2_n3), .B(Key2[26]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[26]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_6_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[26]), .ZN(
        prince_rounds_AddKey2_XORInst_6_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_6_3_U2 ( .A(
        prince_rounds_AddKey2_XORInst_6_3_n3), .B(Key2[27]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[27]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_6_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[27]), .ZN(
        prince_rounds_AddKey2_XORInst_6_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_7_0_U2 ( .A(
        prince_rounds_AddKey2_XORInst_7_0_n3), .B(Key2[28]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[28]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_7_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[28]), .ZN(
        prince_rounds_AddKey2_XORInst_7_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_7_1_U2 ( .A(
        prince_rounds_AddKey2_XORInst_7_1_n3), .B(Key2[29]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[29]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_7_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[29]), .ZN(
        prince_rounds_AddKey2_XORInst_7_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_7_2_U2 ( .A(
        prince_rounds_AddKey2_XORInst_7_2_n3), .B(Key2[30]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[30]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_7_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[30]), .ZN(
        prince_rounds_AddKey2_XORInst_7_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_7_3_U2 ( .A(
        prince_rounds_AddKey2_XORInst_7_3_n3), .B(Key2[31]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[31]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_7_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[31]), .ZN(
        prince_rounds_AddKey2_XORInst_7_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_8_0_U2 ( .A(
        prince_rounds_AddKey2_XORInst_8_0_n3), .B(Key2[32]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[32]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_8_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[32]), .ZN(
        prince_rounds_AddKey2_XORInst_8_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_8_1_U2 ( .A(
        prince_rounds_AddKey2_XORInst_8_1_n3), .B(Key2[33]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[33]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_8_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[33]), .ZN(
        prince_rounds_AddKey2_XORInst_8_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_8_2_U2 ( .A(
        prince_rounds_AddKey2_XORInst_8_2_n3), .B(Key2[34]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[34]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_8_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[34]), .ZN(
        prince_rounds_AddKey2_XORInst_8_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_8_3_U2 ( .A(
        prince_rounds_AddKey2_XORInst_8_3_n3), .B(Key2[35]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[35]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_8_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[35]), .ZN(
        prince_rounds_AddKey2_XORInst_8_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_9_0_U2 ( .A(
        prince_rounds_AddKey2_XORInst_9_0_n3), .B(Key2[36]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[36]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_9_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[36]), .ZN(
        prince_rounds_AddKey2_XORInst_9_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_9_1_U2 ( .A(
        prince_rounds_AddKey2_XORInst_9_1_n3), .B(Key2[37]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[37]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_9_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[37]), .ZN(
        prince_rounds_AddKey2_XORInst_9_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_9_2_U2 ( .A(
        prince_rounds_AddKey2_XORInst_9_2_n3), .B(Key2[38]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[38]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_9_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[38]), .ZN(
        prince_rounds_AddKey2_XORInst_9_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_9_3_U2 ( .A(
        prince_rounds_AddKey2_XORInst_9_3_n3), .B(Key2[39]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[39]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_9_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[39]), .ZN(
        prince_rounds_AddKey2_XORInst_9_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_10_0_U2 ( .A(
        prince_rounds_AddKey2_XORInst_10_0_n3), .B(Key2[40]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[40]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_10_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[40]), .ZN(
        prince_rounds_AddKey2_XORInst_10_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_10_1_U2 ( .A(
        prince_rounds_AddKey2_XORInst_10_1_n3), .B(Key2[41]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[41]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_10_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[41]), .ZN(
        prince_rounds_AddKey2_XORInst_10_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_10_2_U2 ( .A(
        prince_rounds_AddKey2_XORInst_10_2_n3), .B(Key2[42]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[42]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_10_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[42]), .ZN(
        prince_rounds_AddKey2_XORInst_10_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_10_3_U2 ( .A(
        prince_rounds_AddKey2_XORInst_10_3_n3), .B(Key2[43]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[43]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_10_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[43]), .ZN(
        prince_rounds_AddKey2_XORInst_10_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_11_0_U2 ( .A(
        prince_rounds_AddKey2_XORInst_11_0_n3), .B(Key2[44]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[44]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_11_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[44]), .ZN(
        prince_rounds_AddKey2_XORInst_11_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_11_1_U2 ( .A(
        prince_rounds_AddKey2_XORInst_11_1_n3), .B(Key2[45]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[45]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_11_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[45]), .ZN(
        prince_rounds_AddKey2_XORInst_11_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_11_2_U2 ( .A(
        prince_rounds_AddKey2_XORInst_11_2_n3), .B(Key2[46]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[46]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_11_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[46]), .ZN(
        prince_rounds_AddKey2_XORInst_11_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_11_3_U2 ( .A(
        prince_rounds_AddKey2_XORInst_11_3_n3), .B(Key2[47]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[47]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_11_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[47]), .ZN(
        prince_rounds_AddKey2_XORInst_11_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_12_0_U2 ( .A(
        prince_rounds_AddKey2_XORInst_12_0_n3), .B(Key2[48]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[48]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_12_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[48]), .ZN(
        prince_rounds_AddKey2_XORInst_12_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_12_1_U2 ( .A(
        prince_rounds_AddKey2_XORInst_12_1_n3), .B(Key2[49]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[49]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_12_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[49]), .ZN(
        prince_rounds_AddKey2_XORInst_12_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_12_2_U2 ( .A(
        prince_rounds_AddKey2_XORInst_12_2_n3), .B(Key2[50]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[50]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_12_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[50]), .ZN(
        prince_rounds_AddKey2_XORInst_12_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_12_3_U2 ( .A(
        prince_rounds_AddKey2_XORInst_12_3_n3), .B(Key2[51]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[51]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_12_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[51]), .ZN(
        prince_rounds_AddKey2_XORInst_12_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_13_0_U2 ( .A(
        prince_rounds_AddKey2_XORInst_13_0_n3), .B(Key2[52]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[52]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_13_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[52]), .ZN(
        prince_rounds_AddKey2_XORInst_13_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_13_1_U2 ( .A(
        prince_rounds_AddKey2_XORInst_13_1_n3), .B(Key2[53]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[53]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_13_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[53]), .ZN(
        prince_rounds_AddKey2_XORInst_13_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_13_2_U2 ( .A(
        prince_rounds_AddKey2_XORInst_13_2_n3), .B(Key2[54]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[54]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_13_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[54]), .ZN(
        prince_rounds_AddKey2_XORInst_13_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_13_3_U2 ( .A(
        prince_rounds_AddKey2_XORInst_13_3_n3), .B(Key2[55]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[55]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_13_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[55]), .ZN(
        prince_rounds_AddKey2_XORInst_13_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_14_0_U2 ( .A(
        prince_rounds_AddKey2_XORInst_14_0_n3), .B(Key2[56]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[56]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_14_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[56]), .ZN(
        prince_rounds_AddKey2_XORInst_14_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_14_1_U2 ( .A(
        prince_rounds_AddKey2_XORInst_14_1_n3), .B(Key2[57]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[57]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_14_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[57]), .ZN(
        prince_rounds_AddKey2_XORInst_14_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_14_2_U2 ( .A(
        prince_rounds_AddKey2_XORInst_14_2_n3), .B(Key2[58]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[58]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_14_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[58]), .ZN(
        prince_rounds_AddKey2_XORInst_14_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_14_3_U2 ( .A(
        prince_rounds_AddKey2_XORInst_14_3_n3), .B(Key2[59]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[59]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_14_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[59]), .ZN(
        prince_rounds_AddKey2_XORInst_14_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_15_0_U2 ( .A(
        prince_rounds_AddKey2_XORInst_15_0_n3), .B(Key2[60]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[60]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_15_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[60]), .ZN(
        prince_rounds_AddKey2_XORInst_15_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_15_1_U2 ( .A(
        prince_rounds_AddKey2_XORInst_15_1_n3), .B(Key2[61]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[61]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_15_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[61]), .ZN(
        prince_rounds_AddKey2_XORInst_15_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_15_2_U2 ( .A(
        prince_rounds_AddKey2_XORInst_15_2_n3), .B(Key2[62]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[62]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_15_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[62]), .ZN(
        prince_rounds_AddKey2_XORInst_15_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_15_3_U2 ( .A(
        prince_rounds_AddKey2_XORInst_15_3_n3), .B(Key2[63]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s2[63]) );
  XNOR2_X1 prince_rounds_AddKey2_XORInst_15_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s2[63]), .ZN(
        prince_rounds_AddKey2_XORInst_15_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_0_0_U2 ( .A(
        prince_rounds_AddKey3_XORInst_0_0_n3), .B(Key3[0]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[0]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_0_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[0]), .ZN(
        prince_rounds_AddKey3_XORInst_0_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_0_1_U2 ( .A(
        prince_rounds_AddKey3_XORInst_0_1_n3), .B(Key3[1]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[1]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_0_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[1]), .ZN(
        prince_rounds_AddKey3_XORInst_0_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_0_2_U2 ( .A(
        prince_rounds_AddKey3_XORInst_0_2_n3), .B(Key3[2]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[2]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_0_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[2]), .ZN(
        prince_rounds_AddKey3_XORInst_0_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_0_3_U2 ( .A(
        prince_rounds_AddKey3_XORInst_0_3_n3), .B(Key3[3]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[3]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_0_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[3]), .ZN(
        prince_rounds_AddKey3_XORInst_0_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_1_0_U2 ( .A(
        prince_rounds_AddKey3_XORInst_1_0_n3), .B(Key3[4]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[4]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_1_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[4]), .ZN(
        prince_rounds_AddKey3_XORInst_1_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_1_1_U2 ( .A(
        prince_rounds_AddKey3_XORInst_1_1_n3), .B(Key3[5]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[5]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_1_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[5]), .ZN(
        prince_rounds_AddKey3_XORInst_1_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_1_2_U2 ( .A(
        prince_rounds_AddKey3_XORInst_1_2_n3), .B(Key3[6]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[6]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_1_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[6]), .ZN(
        prince_rounds_AddKey3_XORInst_1_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_1_3_U2 ( .A(
        prince_rounds_AddKey3_XORInst_1_3_n3), .B(Key3[7]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[7]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_1_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[7]), .ZN(
        prince_rounds_AddKey3_XORInst_1_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_2_0_U2 ( .A(
        prince_rounds_AddKey3_XORInst_2_0_n3), .B(Key3[8]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[8]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_2_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[8]), .ZN(
        prince_rounds_AddKey3_XORInst_2_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_2_1_U2 ( .A(
        prince_rounds_AddKey3_XORInst_2_1_n3), .B(Key3[9]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[9]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_2_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[9]), .ZN(
        prince_rounds_AddKey3_XORInst_2_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_2_2_U2 ( .A(
        prince_rounds_AddKey3_XORInst_2_2_n3), .B(Key3[10]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[10]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_2_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[10]), .ZN(
        prince_rounds_AddKey3_XORInst_2_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_2_3_U2 ( .A(
        prince_rounds_AddKey3_XORInst_2_3_n3), .B(Key3[11]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[11]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_2_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[11]), .ZN(
        prince_rounds_AddKey3_XORInst_2_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_3_0_U2 ( .A(
        prince_rounds_AddKey3_XORInst_3_0_n3), .B(Key3[12]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[12]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_3_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[12]), .ZN(
        prince_rounds_AddKey3_XORInst_3_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_3_1_U2 ( .A(
        prince_rounds_AddKey3_XORInst_3_1_n3), .B(Key3[13]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[13]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_3_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[13]), .ZN(
        prince_rounds_AddKey3_XORInst_3_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_3_2_U2 ( .A(
        prince_rounds_AddKey3_XORInst_3_2_n3), .B(Key3[14]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[14]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_3_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[14]), .ZN(
        prince_rounds_AddKey3_XORInst_3_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_3_3_U2 ( .A(
        prince_rounds_AddKey3_XORInst_3_3_n3), .B(Key3[15]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[15]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_3_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[15]), .ZN(
        prince_rounds_AddKey3_XORInst_3_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_4_0_U2 ( .A(
        prince_rounds_AddKey3_XORInst_4_0_n3), .B(Key3[16]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[16]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_4_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[16]), .ZN(
        prince_rounds_AddKey3_XORInst_4_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_4_1_U2 ( .A(
        prince_rounds_AddKey3_XORInst_4_1_n3), .B(Key3[17]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[17]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_4_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[17]), .ZN(
        prince_rounds_AddKey3_XORInst_4_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_4_2_U2 ( .A(
        prince_rounds_AddKey3_XORInst_4_2_n3), .B(Key3[18]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[18]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_4_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[18]), .ZN(
        prince_rounds_AddKey3_XORInst_4_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_4_3_U2 ( .A(
        prince_rounds_AddKey3_XORInst_4_3_n3), .B(Key3[19]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[19]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_4_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[19]), .ZN(
        prince_rounds_AddKey3_XORInst_4_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_5_0_U2 ( .A(
        prince_rounds_AddKey3_XORInst_5_0_n3), .B(Key3[20]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[20]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_5_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[20]), .ZN(
        prince_rounds_AddKey3_XORInst_5_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_5_1_U2 ( .A(
        prince_rounds_AddKey3_XORInst_5_1_n3), .B(Key3[21]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[21]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_5_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[21]), .ZN(
        prince_rounds_AddKey3_XORInst_5_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_5_2_U2 ( .A(
        prince_rounds_AddKey3_XORInst_5_2_n3), .B(Key3[22]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[22]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_5_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[22]), .ZN(
        prince_rounds_AddKey3_XORInst_5_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_5_3_U2 ( .A(
        prince_rounds_AddKey3_XORInst_5_3_n3), .B(Key3[23]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[23]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_5_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[23]), .ZN(
        prince_rounds_AddKey3_XORInst_5_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_6_0_U2 ( .A(
        prince_rounds_AddKey3_XORInst_6_0_n3), .B(Key3[24]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[24]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_6_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[24]), .ZN(
        prince_rounds_AddKey3_XORInst_6_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_6_1_U2 ( .A(
        prince_rounds_AddKey3_XORInst_6_1_n3), .B(Key3[25]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[25]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_6_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[25]), .ZN(
        prince_rounds_AddKey3_XORInst_6_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_6_2_U2 ( .A(
        prince_rounds_AddKey3_XORInst_6_2_n3), .B(Key3[26]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[26]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_6_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[26]), .ZN(
        prince_rounds_AddKey3_XORInst_6_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_6_3_U2 ( .A(
        prince_rounds_AddKey3_XORInst_6_3_n3), .B(Key3[27]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[27]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_6_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[27]), .ZN(
        prince_rounds_AddKey3_XORInst_6_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_7_0_U2 ( .A(
        prince_rounds_AddKey3_XORInst_7_0_n3), .B(Key3[28]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[28]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_7_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[28]), .ZN(
        prince_rounds_AddKey3_XORInst_7_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_7_1_U2 ( .A(
        prince_rounds_AddKey3_XORInst_7_1_n3), .B(Key3[29]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[29]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_7_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[29]), .ZN(
        prince_rounds_AddKey3_XORInst_7_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_7_2_U2 ( .A(
        prince_rounds_AddKey3_XORInst_7_2_n3), .B(Key3[30]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[30]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_7_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[30]), .ZN(
        prince_rounds_AddKey3_XORInst_7_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_7_3_U2 ( .A(
        prince_rounds_AddKey3_XORInst_7_3_n3), .B(Key3[31]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[31]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_7_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[31]), .ZN(
        prince_rounds_AddKey3_XORInst_7_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_8_0_U2 ( .A(
        prince_rounds_AddKey3_XORInst_8_0_n3), .B(Key3[32]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[32]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_8_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[32]), .ZN(
        prince_rounds_AddKey3_XORInst_8_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_8_1_U2 ( .A(
        prince_rounds_AddKey3_XORInst_8_1_n3), .B(Key3[33]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[33]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_8_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[33]), .ZN(
        prince_rounds_AddKey3_XORInst_8_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_8_2_U2 ( .A(
        prince_rounds_AddKey3_XORInst_8_2_n3), .B(Key3[34]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[34]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_8_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[34]), .ZN(
        prince_rounds_AddKey3_XORInst_8_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_8_3_U2 ( .A(
        prince_rounds_AddKey3_XORInst_8_3_n3), .B(Key3[35]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[35]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_8_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[35]), .ZN(
        prince_rounds_AddKey3_XORInst_8_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_9_0_U2 ( .A(
        prince_rounds_AddKey3_XORInst_9_0_n3), .B(Key3[36]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[36]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_9_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[36]), .ZN(
        prince_rounds_AddKey3_XORInst_9_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_9_1_U2 ( .A(
        prince_rounds_AddKey3_XORInst_9_1_n3), .B(Key3[37]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[37]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_9_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[37]), .ZN(
        prince_rounds_AddKey3_XORInst_9_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_9_2_U2 ( .A(
        prince_rounds_AddKey3_XORInst_9_2_n3), .B(Key3[38]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[38]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_9_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[38]), .ZN(
        prince_rounds_AddKey3_XORInst_9_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_9_3_U2 ( .A(
        prince_rounds_AddKey3_XORInst_9_3_n3), .B(Key3[39]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[39]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_9_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[39]), .ZN(
        prince_rounds_AddKey3_XORInst_9_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_10_0_U2 ( .A(
        prince_rounds_AddKey3_XORInst_10_0_n3), .B(Key3[40]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[40]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_10_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[40]), .ZN(
        prince_rounds_AddKey3_XORInst_10_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_10_1_U2 ( .A(
        prince_rounds_AddKey3_XORInst_10_1_n3), .B(Key3[41]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[41]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_10_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[41]), .ZN(
        prince_rounds_AddKey3_XORInst_10_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_10_2_U2 ( .A(
        prince_rounds_AddKey3_XORInst_10_2_n3), .B(Key3[42]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[42]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_10_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[42]), .ZN(
        prince_rounds_AddKey3_XORInst_10_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_10_3_U2 ( .A(
        prince_rounds_AddKey3_XORInst_10_3_n3), .B(Key3[43]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[43]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_10_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[43]), .ZN(
        prince_rounds_AddKey3_XORInst_10_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_11_0_U2 ( .A(
        prince_rounds_AddKey3_XORInst_11_0_n3), .B(Key3[44]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[44]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_11_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[44]), .ZN(
        prince_rounds_AddKey3_XORInst_11_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_11_1_U2 ( .A(
        prince_rounds_AddKey3_XORInst_11_1_n3), .B(Key3[45]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[45]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_11_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[45]), .ZN(
        prince_rounds_AddKey3_XORInst_11_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_11_2_U2 ( .A(
        prince_rounds_AddKey3_XORInst_11_2_n3), .B(Key3[46]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[46]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_11_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[46]), .ZN(
        prince_rounds_AddKey3_XORInst_11_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_11_3_U2 ( .A(
        prince_rounds_AddKey3_XORInst_11_3_n3), .B(Key3[47]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[47]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_11_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[47]), .ZN(
        prince_rounds_AddKey3_XORInst_11_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_12_0_U2 ( .A(
        prince_rounds_AddKey3_XORInst_12_0_n3), .B(Key3[48]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[48]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_12_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[48]), .ZN(
        prince_rounds_AddKey3_XORInst_12_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_12_1_U2 ( .A(
        prince_rounds_AddKey3_XORInst_12_1_n3), .B(Key3[49]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[49]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_12_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[49]), .ZN(
        prince_rounds_AddKey3_XORInst_12_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_12_2_U2 ( .A(
        prince_rounds_AddKey3_XORInst_12_2_n3), .B(Key3[50]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[50]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_12_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[50]), .ZN(
        prince_rounds_AddKey3_XORInst_12_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_12_3_U2 ( .A(
        prince_rounds_AddKey3_XORInst_12_3_n3), .B(Key3[51]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[51]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_12_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[51]), .ZN(
        prince_rounds_AddKey3_XORInst_12_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_13_0_U2 ( .A(
        prince_rounds_AddKey3_XORInst_13_0_n3), .B(Key3[52]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[52]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_13_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[52]), .ZN(
        prince_rounds_AddKey3_XORInst_13_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_13_1_U2 ( .A(
        prince_rounds_AddKey3_XORInst_13_1_n3), .B(Key3[53]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[53]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_13_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[53]), .ZN(
        prince_rounds_AddKey3_XORInst_13_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_13_2_U2 ( .A(
        prince_rounds_AddKey3_XORInst_13_2_n3), .B(Key3[54]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[54]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_13_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[54]), .ZN(
        prince_rounds_AddKey3_XORInst_13_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_13_3_U2 ( .A(
        prince_rounds_AddKey3_XORInst_13_3_n3), .B(Key3[55]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[55]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_13_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[55]), .ZN(
        prince_rounds_AddKey3_XORInst_13_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_14_0_U2 ( .A(
        prince_rounds_AddKey3_XORInst_14_0_n3), .B(Key3[56]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[56]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_14_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[56]), .ZN(
        prince_rounds_AddKey3_XORInst_14_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_14_1_U2 ( .A(
        prince_rounds_AddKey3_XORInst_14_1_n3), .B(Key3[57]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[57]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_14_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[57]), .ZN(
        prince_rounds_AddKey3_XORInst_14_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_14_2_U2 ( .A(
        prince_rounds_AddKey3_XORInst_14_2_n3), .B(Key3[58]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[58]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_14_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[58]), .ZN(
        prince_rounds_AddKey3_XORInst_14_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_14_3_U2 ( .A(
        prince_rounds_AddKey3_XORInst_14_3_n3), .B(Key3[59]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[59]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_14_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[59]), .ZN(
        prince_rounds_AddKey3_XORInst_14_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_15_0_U2 ( .A(
        prince_rounds_AddKey3_XORInst_15_0_n3), .B(Key3[60]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[60]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_15_0_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[60]), .ZN(
        prince_rounds_AddKey3_XORInst_15_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_15_1_U2 ( .A(
        prince_rounds_AddKey3_XORInst_15_1_n3), .B(Key3[61]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[61]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_15_1_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[61]), .ZN(
        prince_rounds_AddKey3_XORInst_15_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_15_2_U2 ( .A(
        prince_rounds_AddKey3_XORInst_15_2_n3), .B(Key3[62]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[62]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_15_2_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[62]), .ZN(
        prince_rounds_AddKey3_XORInst_15_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_15_3_U2 ( .A(
        prince_rounds_AddKey3_XORInst_15_3_n3), .B(Key3[63]), .ZN(
        prince_rounds_round_inputXORkeyRCON_s3[63]) );
  XNOR2_X1 prince_rounds_AddKey3_XORInst_15_3_U1 ( .A(1'b0), .B(
        prince_rounds_SR_Result_s3[63]), .ZN(
        prince_rounds_AddKey3_XORInst_15_3_n3) );
  BUF_X4 prince_rounds_sub_U2 ( .A(roundHalf_Select_Signal), .Z(
        prince_rounds_sub_n4) );
  BUF_X8 prince_rounds_sub_U1 ( .A(roundHalf_Select_Signal), .Z(
        prince_rounds_sub_n3) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s1_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[3]), .B(
        prince_rounds_SR_Result_s1[50]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s1_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[0]), .B(
        prince_rounds_SR_Result_s1[49]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s1_n21), .B(
        prince_rounds_SR_Result_s1[48]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s1_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s1_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s1_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[3]), .B(
        prince_rounds_round_inputXORkeyRCON_s1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s1_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[2]), .B(
        prince_rounds_SR_Result_s1[51]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_InAffin_s1_3_) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_U8 ( .B1(
        prince_rounds_sub_n4), .B2(prince_rounds_round_inputXORkeyRCON_s2[2]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_InAffin_s2_3_) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_U7 ( .A1(
        prince_rounds_sub_n4), .A2(prince_rounds_SR_Result_s2[51]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[3]), .B(
        prince_rounds_SR_Result_s2[50]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2[2]) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_U5 ( .B1(
        prince_rounds_sub_n4), .B2(prince_rounds_round_inputXORkeyRCON_s2[0]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_U4 ( .A1(
        prince_rounds_sub_n4), .A2(prince_rounds_SR_Result_s2[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_n16), .B(
        prince_rounds_SR_Result_s2[48]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_n16) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[3]), .B(
        prince_rounds_round_inputXORkeyRCON_s2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s2_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s3_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[3]), .B(
        prince_rounds_SR_Result_s3[50]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s3_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[0]), .B(
        prince_rounds_SR_Result_s3[49]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s3_n21), .B(
        prince_rounds_SR_Result_s3[48]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s3_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s3[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s3_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s3_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[3]), .B(
        prince_rounds_round_inputXORkeyRCON_s3[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s3_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_Pass_inst_s3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[2]), .B(
        prince_rounds_SR_Result_s3[51]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_InAffin_s3_3_) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[3]), .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_InAffin_s1_3_), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_InAffin_s2_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_InAffin_s3_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_n1), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_n1), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[2]), .B(
        r[36]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_n1)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[3]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3[0]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_1__CF_Inst_U1 ( 
        .A(r[0]), .B(r[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_2__CF_Inst_U1 ( 
        .A(r[1]), .B(r[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_4__CF_Inst_U1 ( 
        .A(r[2]), .B(r[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_5__CF_Inst_U1 ( 
        .A(r[3]), .B(r[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_7__CF_Inst_U1 ( 
        .A(r[4]), .B(r[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_8__CF_Inst_U1 ( 
        .A(r[5]), .B(r[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_11__CF_Inst_U1 ( 
        .A(r[7]), .B(r[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_14__CF_Inst_U1 ( 
        .A(r[9]), .B(r[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_16__CF_Inst_U1 ( 
        .A(r[10]), .B(r[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_17__CF_Inst_U1 ( 
        .A(r[11]), .B(r[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_1_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_1_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst1_InstXOR_1__Compression3_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_1_out1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1[2]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_1_out1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[2]), .B(r[37]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_2_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_2_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_2_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_1__CF_Inst_U1 ( 
        .A(r[12]), .B(r[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_2__CF_Inst_U1 ( 
        .A(r[13]), .B(r[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_4__CF_Inst_U1 ( 
        .A(r[14]), .B(r[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_5__CF_Inst_U1 ( 
        .A(r[15]), .B(r[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_7__CF_Inst_U1 ( 
        .A(r[16]), .B(r[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_8__CF_Inst_U1 ( 
        .A(r[17]), .B(r[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_10__CF_Inst_U1 ( 
        .A(r[18]), .B(r[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_11__CF_Inst_U1 ( 
        .A(r[19]), .B(r[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_13__CF_Inst_U1 ( 
        .A(r[20]), .B(r[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_14__CF_Inst_U1 ( 
        .A(r[21]), .B(r[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_16__CF_Inst_U1 ( 
        .A(r[22]), .B(r[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_17__CF_Inst_U1 ( 
        .A(r[23]), .B(r[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_2_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_2_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_2_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst2_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_2_out1[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_2_out1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2Affine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_2_out2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2Affine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_2_out2[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2Affine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_2_out3[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2Affine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_2_out3[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[2]), .B(1'b0), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s1[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s2[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s3[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_1__CF_Inst_U1 ( 
        .A(r[24]), .B(r[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_2__CF_Inst_U1 ( 
        .A(r[25]), .B(r[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_4__CF_Inst_U1 ( 
        .A(r[26]), .B(r[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_5__CF_Inst_U1 ( 
        .A(r[27]), .B(r[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_7__CF_Inst_U1 ( 
        .A(r[28]), .B(r[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_8__CF_Inst_U1 ( 
        .A(r[29]), .B(r[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_10__CF_Inst_U1 ( 
        .A(r[30]), .B(r[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_11__CF_Inst_U1 ( 
        .A(r[31]), .B(r[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_13__CF_Inst_U1 ( 
        .A(r[32]), .B(r[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_14__CF_Inst_U1 ( 
        .A(r[33]), .B(r[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_16__CF_Inst_U1 ( 
        .A(r[34]), .B(r[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_17__CF_Inst_U1 ( 
        .A(r[35]), .B(r[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_inst3_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_OutputAffine1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out1[3]), .Z(
        prince_rounds_sub_Result_s1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_OutputAffine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out1[0]), .B(
        prince_rounds_sub_Result_s1[2]), .ZN(
        prince_rounds_sub_Inv_Result_s1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_OutputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out1[0]), .Z(
        prince_rounds_sub_Result_s1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_OutputAffine2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out2[3]), .Z(
        prince_rounds_sub_Result_s2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_OutputAffine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out2[0]), .B(
        prince_rounds_sub_Result_s2[2]), .Z(prince_rounds_sub_Inv_Result_s2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_OutputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out2[0]), .Z(
        prince_rounds_sub_Result_s2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_OutputAffine3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out3[3]), .Z(
        prince_rounds_sub_Inv_Result_s3[2]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_OutputAffine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out3[0]), .B(
        prince_rounds_sub_Result_s3[2]), .Z(prince_rounds_sub_Inv_Result_s3[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_OutputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_0_Sub_Q294_3_out3[0]), .Z(
        prince_rounds_sub_Inv_Result_s3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s1_n3), .B(
        prince_rounds_sub_Result_s1[2]), .ZN(prince_rounds_sub_Result_s1[0])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s1_U1 ( .A(
        prince_rounds_sub_Result_s1[1]), .B(prince_rounds_sub_Inv_Result_s1[1]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s2_n3), .B(
        prince_rounds_sub_Result_s2[2]), .ZN(prince_rounds_sub_Result_s2[0])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s2_U1 ( .A(
        prince_rounds_sub_Result_s2[1]), .B(prince_rounds_sub_Inv_Result_s2[1]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s2_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s3_U4 ( .A(
        prince_rounds_sub_Inv_Result_s3[2]), .ZN(
        prince_rounds_sub_Result_s3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s3_n5), .B(
        prince_rounds_sub_Result_s3[1]), .ZN(prince_rounds_sub_Result_s3[0])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s3_U2 ( .A(
        prince_rounds_sub_Result_s3[2]), .B(prince_rounds_sub_Inv_Result_s3[1]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s3_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_0_A_inst_s3_U1 ( .A(
        prince_rounds_sub_Inv_Result_s3[0]), .ZN(
        prince_rounds_sub_Result_s3[1]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s1_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[7]), .B(
        prince_rounds_SR_Result_s1[38]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s1_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[4]), .B(
        prince_rounds_SR_Result_s1[37]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s1_n21), .B(
        prince_rounds_SR_Result_s1[36]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s1_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s1[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s1_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s1_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[7]), .B(
        prince_rounds_round_inputXORkeyRCON_s1[4]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s1_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[6]), .B(
        prince_rounds_SR_Result_s1[39]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_InAffin_s1_3_) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_U8 ( .B1(
        prince_rounds_sub_n4), .B2(prince_rounds_round_inputXORkeyRCON_s2[6]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_InAffin_s2_3_) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_U7 ( .A1(
        prince_rounds_sub_n4), .A2(prince_rounds_SR_Result_s2[39]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[7]), .B(
        prince_rounds_SR_Result_s2[38]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2[2]) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_U5 ( .B1(
        prince_rounds_sub_n4), .B2(prince_rounds_round_inputXORkeyRCON_s2[4]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_U4 ( .A1(
        prince_rounds_sub_n4), .A2(prince_rounds_SR_Result_s2[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_n16), .B(
        prince_rounds_SR_Result_s2[36]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[5]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_n16) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[7]), .B(
        prince_rounds_round_inputXORkeyRCON_s2[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s2_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s3_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[7]), .B(
        prince_rounds_SR_Result_s3[38]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s3_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[4]), .B(
        prince_rounds_SR_Result_s3[37]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s3_n21), .B(
        prince_rounds_SR_Result_s3[36]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s3_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s3[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s3_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s3_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[7]), .B(
        prince_rounds_round_inputXORkeyRCON_s3[4]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s3_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_Pass_inst_s3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[6]), .B(
        prince_rounds_SR_Result_s3[39]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_InAffin_s3_3_) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[3]), .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_InAffin_s1_3_), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_InAffin_s2_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_InAffin_s3_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[2]), .B(
        r[36]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_n3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[3]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3[0]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_1__CF_Inst_U1 ( 
        .A(r[0]), .B(r[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_2__CF_Inst_U1 ( 
        .A(r[1]), .B(r[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_4__CF_Inst_U1 ( 
        .A(r[2]), .B(r[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_5__CF_Inst_U1 ( 
        .A(r[3]), .B(r[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_7__CF_Inst_U1 ( 
        .A(r[4]), .B(r[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_8__CF_Inst_U1 ( 
        .A(r[5]), .B(r[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_11__CF_Inst_U1 ( 
        .A(r[7]), .B(r[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_14__CF_Inst_U1 ( 
        .A(r[9]), .B(r[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_16__CF_Inst_U1 ( 
        .A(r[10]), .B(r[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_17__CF_Inst_U1 ( 
        .A(r[11]), .B(r[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_1_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_1_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst1_InstXOR_1__Compression3_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_1_out1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1[2]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_1_out1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[2]), .B(r[37]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_2_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_2_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_2_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_1__CF_Inst_U1 ( 
        .A(r[12]), .B(r[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_2__CF_Inst_U1 ( 
        .A(r[13]), .B(r[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_4__CF_Inst_U1 ( 
        .A(r[14]), .B(r[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_5__CF_Inst_U1 ( 
        .A(r[15]), .B(r[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_7__CF_Inst_U1 ( 
        .A(r[16]), .B(r[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_8__CF_Inst_U1 ( 
        .A(r[17]), .B(r[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_10__CF_Inst_U1 ( 
        .A(r[18]), .B(r[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_11__CF_Inst_U1 ( 
        .A(r[19]), .B(r[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_13__CF_Inst_U1 ( 
        .A(r[20]), .B(r[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_14__CF_Inst_U1 ( 
        .A(r[21]), .B(r[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_16__CF_Inst_U1 ( 
        .A(r[22]), .B(r[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_17__CF_Inst_U1 ( 
        .A(r[23]), .B(r[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_2_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_2_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_2_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst2_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_2_out1[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_2_out1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2Affine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_2_out2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2Affine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_2_out2[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2Affine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_2_out3[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2Affine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_2_out3[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[2]), .B(1'b0), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s1[6]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s2[6]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s3[6]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_1__CF_Inst_U1 ( 
        .A(r[24]), .B(r[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_2__CF_Inst_U1 ( 
        .A(r[25]), .B(r[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_4__CF_Inst_U1 ( 
        .A(r[26]), .B(r[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_5__CF_Inst_U1 ( 
        .A(r[27]), .B(r[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_7__CF_Inst_U1 ( 
        .A(r[28]), .B(r[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_8__CF_Inst_U1 ( 
        .A(r[29]), .B(r[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_10__CF_Inst_U1 ( 
        .A(r[30]), .B(r[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_11__CF_Inst_U1 ( 
        .A(r[31]), .B(r[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_13__CF_Inst_U1 ( 
        .A(r[32]), .B(r[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_14__CF_Inst_U1 ( 
        .A(r[33]), .B(r[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_16__CF_Inst_U1 ( 
        .A(r[34]), .B(r[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_17__CF_Inst_U1 ( 
        .A(r[35]), .B(r[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_inst3_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_OutputAffine1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out1[3]), .Z(
        prince_rounds_sub_Result_s1[7]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_OutputAffine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out1[0]), .B(
        prince_rounds_sub_Result_s1[6]), .ZN(
        prince_rounds_sub_Inv_Result_s1[5]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_OutputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out1[0]), .Z(
        prince_rounds_sub_Result_s1[5]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_OutputAffine2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out2[3]), .Z(
        prince_rounds_sub_Result_s2[7]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_OutputAffine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out2[0]), .B(
        prince_rounds_sub_Result_s2[6]), .Z(prince_rounds_sub_Inv_Result_s2[5]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_OutputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out2[0]), .Z(
        prince_rounds_sub_Result_s2[5]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_OutputAffine3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out3[3]), .Z(
        prince_rounds_sub_Inv_Result_s3[6]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_OutputAffine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out3[0]), .B(
        prince_rounds_sub_Result_s3[6]), .Z(prince_rounds_sub_Inv_Result_s3[5]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_OutputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_1_Sub_Q294_3_out3[0]), .Z(
        prince_rounds_sub_Inv_Result_s3[4]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s1_n3), .B(
        prince_rounds_sub_Result_s1[6]), .ZN(prince_rounds_sub_Result_s1[4])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s1_U1 ( .A(
        prince_rounds_sub_Result_s1[5]), .B(prince_rounds_sub_Inv_Result_s1[5]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s2_n3), .B(
        prince_rounds_sub_Result_s2[6]), .ZN(prince_rounds_sub_Result_s2[4])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s2_U1 ( .A(
        prince_rounds_sub_Result_s2[5]), .B(prince_rounds_sub_Inv_Result_s2[5]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s2_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s3_U4 ( .A(
        prince_rounds_sub_Inv_Result_s3[6]), .ZN(
        prince_rounds_sub_Result_s3[7]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s3_n5), .B(
        prince_rounds_sub_Result_s3[5]), .ZN(prince_rounds_sub_Result_s3[4])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s3_U2 ( .A(
        prince_rounds_sub_Result_s3[6]), .B(prince_rounds_sub_Inv_Result_s3[5]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s3_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_1_A_inst_s3_U1 ( .A(
        prince_rounds_sub_Inv_Result_s3[4]), .ZN(
        prince_rounds_sub_Result_s3[5]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s1_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[11]), .B(
        prince_rounds_SR_Result_s1[26]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s1_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[8]), .B(
        prince_rounds_SR_Result_s1[25]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s1_n21), .B(
        prince_rounds_SR_Result_s1[24]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s1_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s1[9]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s1_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s1_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[11]), .B(
        prince_rounds_round_inputXORkeyRCON_s1[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s1_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[10]), .B(
        prince_rounds_SR_Result_s1[27]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_InAffin_s1_3_) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_U8 ( .B1(
        prince_rounds_sub_n4), .B2(prince_rounds_round_inputXORkeyRCON_s2[10]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_InAffin_s2_3_) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_U7 ( .A1(
        prince_rounds_sub_n4), .A2(prince_rounds_SR_Result_s2[27]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[11]), .B(
        prince_rounds_SR_Result_s2[26]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2[2]) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_U5 ( .B1(
        prince_rounds_sub_n4), .B2(prince_rounds_round_inputXORkeyRCON_s2[8]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_U4 ( .A1(
        prince_rounds_sub_n4), .A2(prince_rounds_SR_Result_s2[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_n16), .B(
        prince_rounds_SR_Result_s2[24]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[9]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_n16) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[11]), .B(
        prince_rounds_round_inputXORkeyRCON_s2[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s2_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s3_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[11]), .B(
        prince_rounds_SR_Result_s3[26]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s3_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[8]), .B(
        prince_rounds_SR_Result_s3[25]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s3_n21), .B(
        prince_rounds_SR_Result_s3[24]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s3_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s3[9]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s3_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s3_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[11]), .B(
        prince_rounds_round_inputXORkeyRCON_s3[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s3_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_Pass_inst_s3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[10]), .B(
        prince_rounds_SR_Result_s3[27]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_InAffin_s3_3_) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[3]), .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_InAffin_s1_3_), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_InAffin_s2_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_InAffin_s3_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[2]), .B(
        r[36]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_n3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[3]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3[0]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_1__CF_Inst_U1 ( 
        .A(r[0]), .B(r[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_2__CF_Inst_U1 ( 
        .A(r[1]), .B(r[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_4__CF_Inst_U1 ( 
        .A(r[2]), .B(r[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_5__CF_Inst_U1 ( 
        .A(r[3]), .B(r[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_7__CF_Inst_U1 ( 
        .A(r[4]), .B(r[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_8__CF_Inst_U1 ( 
        .A(r[5]), .B(r[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_11__CF_Inst_U1 ( 
        .A(r[7]), .B(r[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_14__CF_Inst_U1 ( 
        .A(r[9]), .B(r[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_16__CF_Inst_U1 ( 
        .A(r[10]), .B(r[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_17__CF_Inst_U1 ( 
        .A(r[11]), .B(r[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_1_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_1_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst1_InstXOR_1__Compression3_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_1_out1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1[2]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_1_out1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[2]), .B(r[37]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_2_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_2_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_2_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_1__CF_Inst_U1 ( 
        .A(r[12]), .B(r[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_2__CF_Inst_U1 ( 
        .A(r[13]), .B(r[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_4__CF_Inst_U1 ( 
        .A(r[14]), .B(r[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_5__CF_Inst_U1 ( 
        .A(r[15]), .B(r[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_7__CF_Inst_U1 ( 
        .A(r[16]), .B(r[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_8__CF_Inst_U1 ( 
        .A(r[17]), .B(r[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_10__CF_Inst_U1 ( 
        .A(r[18]), .B(r[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_11__CF_Inst_U1 ( 
        .A(r[19]), .B(r[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_13__CF_Inst_U1 ( 
        .A(r[20]), .B(r[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_14__CF_Inst_U1 ( 
        .A(r[21]), .B(r[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_16__CF_Inst_U1 ( 
        .A(r[22]), .B(r[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_17__CF_Inst_U1 ( 
        .A(r[23]), .B(r[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_2_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_2_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_2_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst2_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_2_out1[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_2_out1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2Affine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_2_out2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2Affine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_2_out2[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2Affine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_2_out3[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2Affine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_2_out3[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[2]), .B(1'b0), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s1[10]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s2[10]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s3[10]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_1__CF_Inst_U1 ( 
        .A(r[24]), .B(r[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_2__CF_Inst_U1 ( 
        .A(r[25]), .B(r[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_4__CF_Inst_U1 ( 
        .A(r[26]), .B(r[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_5__CF_Inst_U1 ( 
        .A(r[27]), .B(r[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_7__CF_Inst_U1 ( 
        .A(r[28]), .B(r[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_8__CF_Inst_U1 ( 
        .A(r[29]), .B(r[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_10__CF_Inst_U1 ( 
        .A(r[30]), .B(r[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_11__CF_Inst_U1 ( 
        .A(r[31]), .B(r[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_13__CF_Inst_U1 ( 
        .A(r[32]), .B(r[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_14__CF_Inst_U1 ( 
        .A(r[33]), .B(r[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_16__CF_Inst_U1 ( 
        .A(r[34]), .B(r[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_17__CF_Inst_U1 ( 
        .A(r[35]), .B(r[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_inst3_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_OutputAffine1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out1[3]), .Z(
        prince_rounds_sub_Result_s1[11]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_OutputAffine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out1[0]), .B(
        prince_rounds_sub_Result_s1[10]), .ZN(
        prince_rounds_sub_Inv_Result_s1[9]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_OutputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out1[0]), .Z(
        prince_rounds_sub_Result_s1[9]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_OutputAffine2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out2[3]), .Z(
        prince_rounds_sub_Result_s2[11]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_OutputAffine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out2[0]), .B(
        prince_rounds_sub_Result_s2[10]), .Z(
        prince_rounds_sub_Inv_Result_s2[9]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_OutputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out2[0]), .Z(
        prince_rounds_sub_Result_s2[9]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_OutputAffine3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out3[3]), .Z(
        prince_rounds_sub_Inv_Result_s3[10]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_OutputAffine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out3[0]), .B(
        prince_rounds_sub_Result_s3[10]), .Z(
        prince_rounds_sub_Inv_Result_s3[9]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_OutputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_2_Sub_Q294_3_out3[0]), .Z(
        prince_rounds_sub_Inv_Result_s3[8]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s1_n3), .B(
        prince_rounds_sub_Result_s1[10]), .ZN(prince_rounds_sub_Result_s1[8])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s1_U1 ( .A(
        prince_rounds_sub_Result_s1[9]), .B(prince_rounds_sub_Inv_Result_s1[9]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s2_n3), .B(
        prince_rounds_sub_Result_s2[10]), .ZN(prince_rounds_sub_Result_s2[8])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s2_U1 ( .A(
        prince_rounds_sub_Result_s2[9]), .B(prince_rounds_sub_Inv_Result_s2[9]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s2_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s3_U4 ( .A(
        prince_rounds_sub_Inv_Result_s3[10]), .ZN(
        prince_rounds_sub_Result_s3[11]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s3_n5), .B(
        prince_rounds_sub_Result_s3[9]), .ZN(prince_rounds_sub_Result_s3[8])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s3_U2 ( .A(
        prince_rounds_sub_Result_s3[10]), .B(
        prince_rounds_sub_Inv_Result_s3[9]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s3_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_2_A_inst_s3_U1 ( .A(
        prince_rounds_sub_Inv_Result_s3[8]), .ZN(
        prince_rounds_sub_Result_s3[9]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s1_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[15]), .B(
        prince_rounds_SR_Result_s1[14]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s1_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[12]), .B(
        prince_rounds_SR_Result_s1[13]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s1_n21), .B(
        prince_rounds_SR_Result_s1[12]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s1_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s1[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s1_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s1_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[15]), .B(
        prince_rounds_round_inputXORkeyRCON_s1[12]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s1_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[14]), .B(
        prince_rounds_SR_Result_s1[15]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_InAffin_s1_3_) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_U8 ( .B1(
        prince_rounds_sub_n4), .B2(prince_rounds_round_inputXORkeyRCON_s2[14]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_InAffin_s2_3_) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_U7 ( .A1(
        prince_rounds_sub_n4), .A2(prince_rounds_SR_Result_s2[15]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[15]), .B(
        prince_rounds_SR_Result_s2[14]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2[2]) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_U5 ( .B1(
        prince_rounds_sub_n4), .B2(prince_rounds_round_inputXORkeyRCON_s2[12]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_U4 ( .A1(
        prince_rounds_sub_n4), .A2(prince_rounds_SR_Result_s2[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_n16), .B(
        prince_rounds_SR_Result_s2[12]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[13]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_n16) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[15]), .B(
        prince_rounds_round_inputXORkeyRCON_s2[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s2_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s3_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[15]), .B(
        prince_rounds_SR_Result_s3[14]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s3_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[12]), .B(
        prince_rounds_SR_Result_s3[13]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s3_n21), .B(
        prince_rounds_SR_Result_s3[12]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s3_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s3[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s3_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s3_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[15]), .B(
        prince_rounds_round_inputXORkeyRCON_s3[12]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s3_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_Pass_inst_s3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[14]), .B(
        prince_rounds_SR_Result_s3[15]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_InAffin_s3_3_) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[3]), .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_InAffin_s1_3_), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_InAffin_s2_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_InAffin_s3_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[2]), .B(
        r[36]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_n3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[3]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3[0]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_1__CF_Inst_U1 ( 
        .A(r[0]), .B(r[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_2__CF_Inst_U1 ( 
        .A(r[1]), .B(r[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_4__CF_Inst_U1 ( 
        .A(r[2]), .B(r[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_5__CF_Inst_U1 ( 
        .A(r[3]), .B(r[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_7__CF_Inst_U1 ( 
        .A(r[4]), .B(r[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_8__CF_Inst_U1 ( 
        .A(r[5]), .B(r[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_11__CF_Inst_U1 ( 
        .A(r[7]), .B(r[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_14__CF_Inst_U1 ( 
        .A(r[9]), .B(r[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_16__CF_Inst_U1 ( 
        .A(r[10]), .B(r[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_17__CF_Inst_U1 ( 
        .A(r[11]), .B(r[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_1_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_1_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst1_InstXOR_1__Compression3_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_1_out1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1[2]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_1_out1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[2]), .B(r[37]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_2_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_2_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_2_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_1__CF_Inst_U1 ( 
        .A(r[12]), .B(r[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_2__CF_Inst_U1 ( 
        .A(r[13]), .B(r[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_4__CF_Inst_U1 ( 
        .A(r[14]), .B(r[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_5__CF_Inst_U1 ( 
        .A(r[15]), .B(r[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_7__CF_Inst_U1 ( 
        .A(r[16]), .B(r[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_8__CF_Inst_U1 ( 
        .A(r[17]), .B(r[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_10__CF_Inst_U1 ( 
        .A(r[18]), .B(r[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_11__CF_Inst_U1 ( 
        .A(r[19]), .B(r[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_13__CF_Inst_U1 ( 
        .A(r[20]), .B(r[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_14__CF_Inst_U1 ( 
        .A(r[21]), .B(r[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_16__CF_Inst_U1 ( 
        .A(r[22]), .B(r[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_17__CF_Inst_U1 ( 
        .A(r[23]), .B(r[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_2_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_2_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_2_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst2_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_2_out1[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_2_out1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2Affine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_2_out2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2Affine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_2_out2[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2Affine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_2_out3[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2Affine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_2_out3[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[2]), .B(1'b0), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s1[14]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s2[14]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s3[14]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_1__CF_Inst_U1 ( 
        .A(r[24]), .B(r[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_2__CF_Inst_U1 ( 
        .A(r[25]), .B(r[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_4__CF_Inst_U1 ( 
        .A(r[26]), .B(r[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_5__CF_Inst_U1 ( 
        .A(r[27]), .B(r[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_7__CF_Inst_U1 ( 
        .A(r[28]), .B(r[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_8__CF_Inst_U1 ( 
        .A(r[29]), .B(r[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_10__CF_Inst_U1 ( 
        .A(r[30]), .B(r[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_11__CF_Inst_U1 ( 
        .A(r[31]), .B(r[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_13__CF_Inst_U1 ( 
        .A(r[32]), .B(r[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_14__CF_Inst_U1 ( 
        .A(r[33]), .B(r[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_16__CF_Inst_U1 ( 
        .A(r[34]), .B(r[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_17__CF_Inst_U1 ( 
        .A(r[35]), .B(r[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_inst3_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_OutputAffine1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out1[3]), .Z(
        prince_rounds_sub_Result_s1[15]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_OutputAffine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out1[0]), .B(
        prince_rounds_sub_Result_s1[14]), .ZN(
        prince_rounds_sub_Inv_Result_s1[13]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_OutputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out1[0]), .Z(
        prince_rounds_sub_Result_s1[13]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_OutputAffine2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out2[3]), .Z(
        prince_rounds_sub_Result_s2[15]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_OutputAffine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out2[0]), .B(
        prince_rounds_sub_Result_s2[14]), .Z(
        prince_rounds_sub_Inv_Result_s2[13]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_OutputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out2[0]), .Z(
        prince_rounds_sub_Result_s2[13]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_OutputAffine3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out3[3]), .Z(
        prince_rounds_sub_Inv_Result_s3[14]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_OutputAffine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out3[0]), .B(
        prince_rounds_sub_Result_s3[14]), .Z(
        prince_rounds_sub_Inv_Result_s3[13]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_OutputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_3_Sub_Q294_3_out3[0]), .Z(
        prince_rounds_sub_Inv_Result_s3[12]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s1_n3), .B(
        prince_rounds_sub_Result_s1[14]), .ZN(prince_rounds_sub_Result_s1[12])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s1_U1 ( .A(
        prince_rounds_sub_Result_s1[13]), .B(
        prince_rounds_sub_Inv_Result_s1[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s2_n3), .B(
        prince_rounds_sub_Result_s2[14]), .ZN(prince_rounds_sub_Result_s2[12])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s2_U1 ( .A(
        prince_rounds_sub_Result_s2[13]), .B(
        prince_rounds_sub_Inv_Result_s2[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s2_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s3_U4 ( .A(
        prince_rounds_sub_Inv_Result_s3[14]), .ZN(
        prince_rounds_sub_Result_s3[15]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s3_n5), .B(
        prince_rounds_sub_Result_s3[13]), .ZN(prince_rounds_sub_Result_s3[12])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s3_U2 ( .A(
        prince_rounds_sub_Result_s3[14]), .B(
        prince_rounds_sub_Inv_Result_s3[13]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s3_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_3_A_inst_s3_U1 ( .A(
        prince_rounds_sub_Inv_Result_s3[12]), .ZN(
        prince_rounds_sub_Result_s3[13]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s1_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[19]), .B(
        prince_rounds_SR_Result_s1[2]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s1_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[16]), .B(
        prince_rounds_SR_Result_s1[1]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s1_n21), .B(
        prince_rounds_SR_Result_s1[0]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s1_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s1[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s1_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s1_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[19]), .B(
        prince_rounds_round_inputXORkeyRCON_s1[16]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s1_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[18]), .B(
        prince_rounds_SR_Result_s1[3]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_InAffin_s1_3_) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_U8 ( .B1(
        prince_rounds_sub_n4), .B2(prince_rounds_round_inputXORkeyRCON_s2[18]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_InAffin_s2_3_) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_U7 ( .A1(
        prince_rounds_sub_n4), .A2(prince_rounds_SR_Result_s2[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[19]), .B(
        prince_rounds_SR_Result_s2[2]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2[2]) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_U5 ( .B1(
        prince_rounds_sub_n4), .B2(prince_rounds_round_inputXORkeyRCON_s2[16]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_U4 ( .A1(
        prince_rounds_sub_n4), .A2(prince_rounds_SR_Result_s2[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_n16), .B(
        prince_rounds_SR_Result_s2[0]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[17]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_n16) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[19]), .B(
        prince_rounds_round_inputXORkeyRCON_s2[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s2_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s3_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[19]), .B(
        prince_rounds_SR_Result_s3[2]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s3_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[16]), .B(
        prince_rounds_SR_Result_s3[1]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s3_n21), .B(
        prince_rounds_SR_Result_s3[0]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s3_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s3[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s3_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s3_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[19]), .B(
        prince_rounds_round_inputXORkeyRCON_s3[16]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s3_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_Pass_inst_s3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[18]), .B(
        prince_rounds_SR_Result_s3[3]), .S(prince_rounds_sub_n4), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_InAffin_s3_3_) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[3]), .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_InAffin_s1_3_), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_InAffin_s2_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_InAffin_s3_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[2]), .B(
        r[36]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_n3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[3]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3[0]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_1__CF_Inst_U1 ( 
        .A(r[0]), .B(r[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_2__CF_Inst_U1 ( 
        .A(r[1]), .B(r[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_4__CF_Inst_U1 ( 
        .A(r[2]), .B(r[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_5__CF_Inst_U1 ( 
        .A(r[3]), .B(r[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_7__CF_Inst_U1 ( 
        .A(r[4]), .B(r[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_8__CF_Inst_U1 ( 
        .A(r[5]), .B(r[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_11__CF_Inst_U1 ( 
        .A(r[7]), .B(r[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_14__CF_Inst_U1 ( 
        .A(r[9]), .B(r[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_16__CF_Inst_U1 ( 
        .A(r[10]), .B(r[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_17__CF_Inst_U1 ( 
        .A(r[11]), .B(r[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_1_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_1_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst1_InstXOR_1__Compression3_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_1_out1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1[2]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_1_out1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[2]), .B(r[37]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_2_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_2_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_2_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_1__CF_Inst_U1 ( 
        .A(r[12]), .B(r[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_2__CF_Inst_U1 ( 
        .A(r[13]), .B(r[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_4__CF_Inst_U1 ( 
        .A(r[14]), .B(r[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_5__CF_Inst_U1 ( 
        .A(r[15]), .B(r[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_7__CF_Inst_U1 ( 
        .A(r[16]), .B(r[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_8__CF_Inst_U1 ( 
        .A(r[17]), .B(r[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_10__CF_Inst_U1 ( 
        .A(r[18]), .B(r[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_11__CF_Inst_U1 ( 
        .A(r[19]), .B(r[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_13__CF_Inst_U1 ( 
        .A(r[20]), .B(r[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_14__CF_Inst_U1 ( 
        .A(r[21]), .B(r[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_16__CF_Inst_U1 ( 
        .A(r[22]), .B(r[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_17__CF_Inst_U1 ( 
        .A(r[23]), .B(r[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_2_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_2_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_2_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst2_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_2_out1[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_2_out1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2Affine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_2_out2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2Affine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_2_out2[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2Affine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_2_out3[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2Affine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_2_out3[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[2]), .B(1'b0), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s1[18]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s2[18]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s3[18]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_1__CF_Inst_U1 ( 
        .A(r[24]), .B(r[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_2__CF_Inst_U1 ( 
        .A(r[25]), .B(r[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_4__CF_Inst_U1 ( 
        .A(r[26]), .B(r[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_5__CF_Inst_U1 ( 
        .A(r[27]), .B(r[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_7__CF_Inst_U1 ( 
        .A(r[28]), .B(r[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_8__CF_Inst_U1 ( 
        .A(r[29]), .B(r[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_10__CF_Inst_U1 ( 
        .A(r[30]), .B(r[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_11__CF_Inst_U1 ( 
        .A(r[31]), .B(r[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_13__CF_Inst_U1 ( 
        .A(r[32]), .B(r[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_14__CF_Inst_U1 ( 
        .A(r[33]), .B(r[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_16__CF_Inst_U1 ( 
        .A(r[34]), .B(r[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_17__CF_Inst_U1 ( 
        .A(r[35]), .B(r[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_inst3_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_OutputAffine1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out1[3]), .Z(
        prince_rounds_sub_Result_s1[19]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_OutputAffine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out1[0]), .B(
        prince_rounds_sub_Result_s1[18]), .ZN(
        prince_rounds_sub_Inv_Result_s1[17]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_OutputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out1[0]), .Z(
        prince_rounds_sub_Result_s1[17]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_OutputAffine2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out2[3]), .Z(
        prince_rounds_sub_Result_s2[19]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_OutputAffine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out2[0]), .B(
        prince_rounds_sub_Result_s2[18]), .Z(
        prince_rounds_sub_Inv_Result_s2[17]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_OutputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out2[0]), .Z(
        prince_rounds_sub_Result_s2[17]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_OutputAffine3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out3[3]), .Z(
        prince_rounds_sub_Inv_Result_s3[18]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_OutputAffine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out3[0]), .B(
        prince_rounds_sub_Result_s3[18]), .Z(
        prince_rounds_sub_Inv_Result_s3[17]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_OutputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_4_Sub_Q294_3_out3[0]), .Z(
        prince_rounds_sub_Inv_Result_s3[16]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s1_n3), .B(
        prince_rounds_sub_Result_s1[18]), .ZN(prince_rounds_sub_Result_s1[16])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s1_U1 ( .A(
        prince_rounds_sub_Result_s1[17]), .B(
        prince_rounds_sub_Inv_Result_s1[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s2_n3), .B(
        prince_rounds_sub_Result_s2[18]), .ZN(prince_rounds_sub_Result_s2[16])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s2_U1 ( .A(
        prince_rounds_sub_Result_s2[17]), .B(
        prince_rounds_sub_Inv_Result_s2[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s2_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s3_U4 ( .A(
        prince_rounds_sub_Inv_Result_s3[18]), .ZN(
        prince_rounds_sub_Result_s3[19]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s3_n5), .B(
        prince_rounds_sub_Result_s3[17]), .ZN(prince_rounds_sub_Result_s3[16])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s3_U2 ( .A(
        prince_rounds_sub_Result_s3[18]), .B(
        prince_rounds_sub_Inv_Result_s3[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s3_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_4_A_inst_s3_U1 ( .A(
        prince_rounds_sub_Inv_Result_s3[16]), .ZN(
        prince_rounds_sub_Result_s3[17]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s1_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[23]), .B(
        prince_rounds_SR_Result_s1[54]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s1_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[20]), .B(
        prince_rounds_SR_Result_s1[53]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s1_n21), .B(
        prince_rounds_SR_Result_s1[52]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s1_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s1[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s1_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s1_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[23]), .B(
        prince_rounds_round_inputXORkeyRCON_s1[20]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s1_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[22]), .B(
        prince_rounds_SR_Result_s1[55]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_InAffin_s1_3_) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_U8 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[22]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_InAffin_s2_3_) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_U7 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[55]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[23]), .B(
        prince_rounds_SR_Result_s2[54]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2[2]) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_U5 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[20]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_U4 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_n16), .B(
        prince_rounds_SR_Result_s2[52]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[21]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_n16) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[23]), .B(
        prince_rounds_round_inputXORkeyRCON_s2[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s2_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s3_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[23]), .B(
        prince_rounds_SR_Result_s3[54]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s3_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[20]), .B(
        prince_rounds_SR_Result_s3[53]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s3_n21), .B(
        prince_rounds_SR_Result_s3[52]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s3_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s3[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s3_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s3_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[23]), .B(
        prince_rounds_round_inputXORkeyRCON_s3[20]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s3_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_Pass_inst_s3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[22]), .B(
        prince_rounds_SR_Result_s3[55]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_InAffin_s3_3_) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[3]), .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_InAffin_s1_3_), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_InAffin_s2_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_InAffin_s3_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[2]), .B(
        r[36]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_n3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[3]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3[0]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_1__CF_Inst_U1 ( 
        .A(r[0]), .B(r[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_2__CF_Inst_U1 ( 
        .A(r[1]), .B(r[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_4__CF_Inst_U1 ( 
        .A(r[2]), .B(r[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_5__CF_Inst_U1 ( 
        .A(r[3]), .B(r[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_7__CF_Inst_U1 ( 
        .A(r[4]), .B(r[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_8__CF_Inst_U1 ( 
        .A(r[5]), .B(r[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_11__CF_Inst_U1 ( 
        .A(r[7]), .B(r[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_14__CF_Inst_U1 ( 
        .A(r[9]), .B(r[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_16__CF_Inst_U1 ( 
        .A(r[10]), .B(r[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_17__CF_Inst_U1 ( 
        .A(r[11]), .B(r[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_1_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_1_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst1_InstXOR_1__Compression3_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_1_out1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1[2]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_1_out1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[2]), .B(r[37]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_2_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_2_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_2_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_1__CF_Inst_U1 ( 
        .A(r[12]), .B(r[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_2__CF_Inst_U1 ( 
        .A(r[13]), .B(r[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_4__CF_Inst_U1 ( 
        .A(r[14]), .B(r[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_5__CF_Inst_U1 ( 
        .A(r[15]), .B(r[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_7__CF_Inst_U1 ( 
        .A(r[16]), .B(r[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_8__CF_Inst_U1 ( 
        .A(r[17]), .B(r[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_10__CF_Inst_U1 ( 
        .A(r[18]), .B(r[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_11__CF_Inst_U1 ( 
        .A(r[19]), .B(r[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_13__CF_Inst_U1 ( 
        .A(r[20]), .B(r[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_14__CF_Inst_U1 ( 
        .A(r[21]), .B(r[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_16__CF_Inst_U1 ( 
        .A(r[22]), .B(r[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_17__CF_Inst_U1 ( 
        .A(r[23]), .B(r[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_2_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_2_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_2_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst2_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_2_out1[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_2_out1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2Affine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_2_out2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2Affine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_2_out2[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2Affine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_2_out3[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2Affine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_2_out3[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[2]), .B(1'b0), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s1[22]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s2[22]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s3[22]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_1__CF_Inst_U1 ( 
        .A(r[24]), .B(r[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_2__CF_Inst_U1 ( 
        .A(r[25]), .B(r[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_4__CF_Inst_U1 ( 
        .A(r[26]), .B(r[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_5__CF_Inst_U1 ( 
        .A(r[27]), .B(r[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_7__CF_Inst_U1 ( 
        .A(r[28]), .B(r[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_8__CF_Inst_U1 ( 
        .A(r[29]), .B(r[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_10__CF_Inst_U1 ( 
        .A(r[30]), .B(r[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_11__CF_Inst_U1 ( 
        .A(r[31]), .B(r[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_13__CF_Inst_U1 ( 
        .A(r[32]), .B(r[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_14__CF_Inst_U1 ( 
        .A(r[33]), .B(r[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_16__CF_Inst_U1 ( 
        .A(r[34]), .B(r[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_17__CF_Inst_U1 ( 
        .A(r[35]), .B(r[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_inst3_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_OutputAffine1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out1[3]), .Z(
        prince_rounds_sub_Result_s1[23]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_OutputAffine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out1[0]), .B(
        prince_rounds_sub_Result_s1[22]), .ZN(
        prince_rounds_sub_Inv_Result_s1[21]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_OutputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out1[0]), .Z(
        prince_rounds_sub_Result_s1[21]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_OutputAffine2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out2[3]), .Z(
        prince_rounds_sub_Result_s2[23]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_OutputAffine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out2[0]), .B(
        prince_rounds_sub_Result_s2[22]), .Z(
        prince_rounds_sub_Inv_Result_s2[21]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_OutputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out2[0]), .Z(
        prince_rounds_sub_Result_s2[21]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_OutputAffine3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out3[3]), .Z(
        prince_rounds_sub_Inv_Result_s3[22]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_OutputAffine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out3[0]), .B(
        prince_rounds_sub_Result_s3[22]), .Z(
        prince_rounds_sub_Inv_Result_s3[21]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_OutputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_5_Sub_Q294_3_out3[0]), .Z(
        prince_rounds_sub_Inv_Result_s3[20]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s1_n3), .B(
        prince_rounds_sub_Result_s1[22]), .ZN(prince_rounds_sub_Result_s1[20])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s1_U1 ( .A(
        prince_rounds_sub_Result_s1[21]), .B(
        prince_rounds_sub_Inv_Result_s1[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s2_n3), .B(
        prince_rounds_sub_Result_s2[22]), .ZN(prince_rounds_sub_Result_s2[20])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s2_U1 ( .A(
        prince_rounds_sub_Result_s2[21]), .B(
        prince_rounds_sub_Inv_Result_s2[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s2_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s3_U4 ( .A(
        prince_rounds_sub_Inv_Result_s3[22]), .ZN(
        prince_rounds_sub_Result_s3[23]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s3_n5), .B(
        prince_rounds_sub_Result_s3[21]), .ZN(prince_rounds_sub_Result_s3[20])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s3_U2 ( .A(
        prince_rounds_sub_Result_s3[22]), .B(
        prince_rounds_sub_Inv_Result_s3[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s3_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_5_A_inst_s3_U1 ( .A(
        prince_rounds_sub_Inv_Result_s3[20]), .ZN(
        prince_rounds_sub_Result_s3[21]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s1_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[27]), .B(
        prince_rounds_SR_Result_s1[42]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s1_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[24]), .B(
        prince_rounds_SR_Result_s1[41]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s1_n21), .B(
        prince_rounds_SR_Result_s1[40]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s1_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s1[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s1_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s1_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[27]), .B(
        prince_rounds_round_inputXORkeyRCON_s1[24]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s1_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[26]), .B(
        prince_rounds_SR_Result_s1[43]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_InAffin_s1_3_) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_U8 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[26]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_InAffin_s2_3_) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_U7 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[43]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[27]), .B(
        prince_rounds_SR_Result_s2[42]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2[2]) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_U5 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[24]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_U4 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_n16), .B(
        prince_rounds_SR_Result_s2[40]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[25]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_n16) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[27]), .B(
        prince_rounds_round_inputXORkeyRCON_s2[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s2_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s3_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[27]), .B(
        prince_rounds_SR_Result_s3[42]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s3_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[24]), .B(
        prince_rounds_SR_Result_s3[41]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s3_n21), .B(
        prince_rounds_SR_Result_s3[40]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s3_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s3[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s3_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s3_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[27]), .B(
        prince_rounds_round_inputXORkeyRCON_s3[24]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s3_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_Pass_inst_s3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[26]), .B(
        prince_rounds_SR_Result_s3[43]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_InAffin_s3_3_) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[3]), .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_InAffin_s1_3_), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_InAffin_s2_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_InAffin_s3_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[2]), .B(
        r[36]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_n3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[3]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3[0]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_1__CF_Inst_U1 ( 
        .A(r[0]), .B(r[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_2__CF_Inst_U1 ( 
        .A(r[1]), .B(r[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_4__CF_Inst_U1 ( 
        .A(r[2]), .B(r[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_5__CF_Inst_U1 ( 
        .A(r[3]), .B(r[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_7__CF_Inst_U1 ( 
        .A(r[4]), .B(r[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_8__CF_Inst_U1 ( 
        .A(r[5]), .B(r[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_11__CF_Inst_U1 ( 
        .A(r[7]), .B(r[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_14__CF_Inst_U1 ( 
        .A(r[9]), .B(r[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_16__CF_Inst_U1 ( 
        .A(r[10]), .B(r[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_17__CF_Inst_U1 ( 
        .A(r[11]), .B(r[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_1_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_1_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst1_InstXOR_1__Compression3_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_1_out1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1[2]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_1_out1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[2]), .B(r[37]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_2_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_2_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_2_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_1__CF_Inst_U1 ( 
        .A(r[12]), .B(r[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_2__CF_Inst_U1 ( 
        .A(r[13]), .B(r[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_4__CF_Inst_U1 ( 
        .A(r[14]), .B(r[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_5__CF_Inst_U1 ( 
        .A(r[15]), .B(r[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_7__CF_Inst_U1 ( 
        .A(r[16]), .B(r[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_8__CF_Inst_U1 ( 
        .A(r[17]), .B(r[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_10__CF_Inst_U1 ( 
        .A(r[18]), .B(r[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_11__CF_Inst_U1 ( 
        .A(r[19]), .B(r[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_13__CF_Inst_U1 ( 
        .A(r[20]), .B(r[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_14__CF_Inst_U1 ( 
        .A(r[21]), .B(r[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_16__CF_Inst_U1 ( 
        .A(r[22]), .B(r[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_17__CF_Inst_U1 ( 
        .A(r[23]), .B(r[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_2_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_2_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_2_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst2_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_2_out1[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_2_out1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2Affine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_2_out2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2Affine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_2_out2[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2Affine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_2_out3[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2Affine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_2_out3[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[2]), .B(1'b0), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s1[26]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s2[26]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s3[26]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_1__CF_Inst_U1 ( 
        .A(r[24]), .B(r[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_2__CF_Inst_U1 ( 
        .A(r[25]), .B(r[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_4__CF_Inst_U1 ( 
        .A(r[26]), .B(r[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_5__CF_Inst_U1 ( 
        .A(r[27]), .B(r[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_7__CF_Inst_U1 ( 
        .A(r[28]), .B(r[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_8__CF_Inst_U1 ( 
        .A(r[29]), .B(r[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_10__CF_Inst_U1 ( 
        .A(r[30]), .B(r[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_11__CF_Inst_U1 ( 
        .A(r[31]), .B(r[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_13__CF_Inst_U1 ( 
        .A(r[32]), .B(r[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_14__CF_Inst_U1 ( 
        .A(r[33]), .B(r[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_16__CF_Inst_U1 ( 
        .A(r[34]), .B(r[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_17__CF_Inst_U1 ( 
        .A(r[35]), .B(r[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_inst3_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_OutputAffine1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out1[3]), .Z(
        prince_rounds_sub_Result_s1[27]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_OutputAffine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out1[0]), .B(
        prince_rounds_sub_Result_s1[26]), .ZN(
        prince_rounds_sub_Inv_Result_s1[25]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_OutputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out1[0]), .Z(
        prince_rounds_sub_Result_s1[25]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_OutputAffine2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out2[3]), .Z(
        prince_rounds_sub_Result_s2[27]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_OutputAffine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out2[0]), .B(
        prince_rounds_sub_Result_s2[26]), .Z(
        prince_rounds_sub_Inv_Result_s2[25]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_OutputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out2[0]), .Z(
        prince_rounds_sub_Result_s2[25]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_OutputAffine3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out3[3]), .Z(
        prince_rounds_sub_Inv_Result_s3[26]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_OutputAffine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out3[0]), .B(
        prince_rounds_sub_Result_s3[26]), .Z(
        prince_rounds_sub_Inv_Result_s3[25]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_OutputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_6_Sub_Q294_3_out3[0]), .Z(
        prince_rounds_sub_Inv_Result_s3[24]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s1_n3), .B(
        prince_rounds_sub_Result_s1[26]), .ZN(prince_rounds_sub_Result_s1[24])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s1_U1 ( .A(
        prince_rounds_sub_Result_s1[25]), .B(
        prince_rounds_sub_Inv_Result_s1[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s2_n3), .B(
        prince_rounds_sub_Result_s2[26]), .ZN(prince_rounds_sub_Result_s2[24])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s2_U1 ( .A(
        prince_rounds_sub_Result_s2[25]), .B(
        prince_rounds_sub_Inv_Result_s2[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s2_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s3_U4 ( .A(
        prince_rounds_sub_Inv_Result_s3[26]), .ZN(
        prince_rounds_sub_Result_s3[27]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s3_n5), .B(
        prince_rounds_sub_Result_s3[25]), .ZN(prince_rounds_sub_Result_s3[24])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s3_U2 ( .A(
        prince_rounds_sub_Result_s3[26]), .B(
        prince_rounds_sub_Inv_Result_s3[25]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s3_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_6_A_inst_s3_U1 ( .A(
        prince_rounds_sub_Inv_Result_s3[24]), .ZN(
        prince_rounds_sub_Result_s3[25]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s1_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[31]), .B(
        prince_rounds_SR_Result_s1[30]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s1_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[28]), .B(
        prince_rounds_SR_Result_s1[29]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s1_n21), .B(
        prince_rounds_SR_Result_s1[28]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s1_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s1[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s1_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s1_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[31]), .B(
        prince_rounds_round_inputXORkeyRCON_s1[28]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s1_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[30]), .B(
        prince_rounds_SR_Result_s1[31]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_InAffin_s1_3_) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_U8 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[30]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_InAffin_s2_3_) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_U7 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[31]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[31]), .B(
        prince_rounds_SR_Result_s2[30]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2[2]) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_U5 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[28]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_U4 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_n16), .B(
        prince_rounds_SR_Result_s2[28]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[29]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_n16) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[31]), .B(
        prince_rounds_round_inputXORkeyRCON_s2[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s2_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s3_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[31]), .B(
        prince_rounds_SR_Result_s3[30]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s3_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[28]), .B(
        prince_rounds_SR_Result_s3[29]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s3_n21), .B(
        prince_rounds_SR_Result_s3[28]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s3_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s3[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s3_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s3_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[31]), .B(
        prince_rounds_round_inputXORkeyRCON_s3[28]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s3_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_Pass_inst_s3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[30]), .B(
        prince_rounds_SR_Result_s3[31]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_InAffin_s3_3_) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[3]), .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_InAffin_s1_3_), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_InAffin_s2_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_InAffin_s3_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[2]), .B(
        r[36]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_n3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[3]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3[0]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_1__CF_Inst_U1 ( 
        .A(r[0]), .B(r[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_2__CF_Inst_U1 ( 
        .A(r[1]), .B(r[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_4__CF_Inst_U1 ( 
        .A(r[2]), .B(r[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_5__CF_Inst_U1 ( 
        .A(r[3]), .B(r[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_7__CF_Inst_U1 ( 
        .A(r[4]), .B(r[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_8__CF_Inst_U1 ( 
        .A(r[5]), .B(r[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_11__CF_Inst_U1 ( 
        .A(r[7]), .B(r[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_14__CF_Inst_U1 ( 
        .A(r[9]), .B(r[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_16__CF_Inst_U1 ( 
        .A(r[10]), .B(r[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_17__CF_Inst_U1 ( 
        .A(r[11]), .B(r[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_1_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_1_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst1_InstXOR_1__Compression3_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_1_out1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1[2]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_1_out1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[2]), .B(r[37]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_2_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_2_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_2_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_1__CF_Inst_U1 ( 
        .A(r[12]), .B(r[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_2__CF_Inst_U1 ( 
        .A(r[13]), .B(r[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_4__CF_Inst_U1 ( 
        .A(r[14]), .B(r[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_5__CF_Inst_U1 ( 
        .A(r[15]), .B(r[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_7__CF_Inst_U1 ( 
        .A(r[16]), .B(r[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_8__CF_Inst_U1 ( 
        .A(r[17]), .B(r[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_10__CF_Inst_U1 ( 
        .A(r[18]), .B(r[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_11__CF_Inst_U1 ( 
        .A(r[19]), .B(r[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_13__CF_Inst_U1 ( 
        .A(r[20]), .B(r[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_14__CF_Inst_U1 ( 
        .A(r[21]), .B(r[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_16__CF_Inst_U1 ( 
        .A(r[22]), .B(r[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_17__CF_Inst_U1 ( 
        .A(r[23]), .B(r[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_2_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_2_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_2_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst2_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_2_out1[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_2_out1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2Affine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_2_out2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2Affine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_2_out2[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2Affine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_2_out3[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2Affine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_2_out3[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[2]), .B(1'b0), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s1[30]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s2[30]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s3[30]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_1__CF_Inst_U1 ( 
        .A(r[24]), .B(r[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_2__CF_Inst_U1 ( 
        .A(r[25]), .B(r[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_4__CF_Inst_U1 ( 
        .A(r[26]), .B(r[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_5__CF_Inst_U1 ( 
        .A(r[27]), .B(r[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_7__CF_Inst_U1 ( 
        .A(r[28]), .B(r[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_8__CF_Inst_U1 ( 
        .A(r[29]), .B(r[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_10__CF_Inst_U1 ( 
        .A(r[30]), .B(r[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_11__CF_Inst_U1 ( 
        .A(r[31]), .B(r[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_13__CF_Inst_U1 ( 
        .A(r[32]), .B(r[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_14__CF_Inst_U1 ( 
        .A(r[33]), .B(r[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_16__CF_Inst_U1 ( 
        .A(r[34]), .B(r[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_17__CF_Inst_U1 ( 
        .A(r[35]), .B(r[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_inst3_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_OutputAffine1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out1[3]), .Z(
        prince_rounds_sub_Result_s1[31]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_OutputAffine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out1[0]), .B(
        prince_rounds_sub_Result_s1[30]), .ZN(
        prince_rounds_sub_Inv_Result_s1[29]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_OutputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out1[0]), .Z(
        prince_rounds_sub_Result_s1[29]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_OutputAffine2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out2[3]), .Z(
        prince_rounds_sub_Result_s2[31]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_OutputAffine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out2[0]), .B(
        prince_rounds_sub_Result_s2[30]), .Z(
        prince_rounds_sub_Inv_Result_s2[29]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_OutputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out2[0]), .Z(
        prince_rounds_sub_Result_s2[29]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_OutputAffine3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out3[3]), .Z(
        prince_rounds_sub_Inv_Result_s3[30]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_OutputAffine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out3[0]), .B(
        prince_rounds_sub_Result_s3[30]), .Z(
        prince_rounds_sub_Inv_Result_s3[29]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_OutputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_7_Sub_Q294_3_out3[0]), .Z(
        prince_rounds_sub_Inv_Result_s3[28]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s1_n3), .B(
        prince_rounds_sub_Result_s1[30]), .ZN(prince_rounds_sub_Result_s1[28])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s1_U1 ( .A(
        prince_rounds_sub_Result_s1[29]), .B(
        prince_rounds_sub_Inv_Result_s1[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s2_n3), .B(
        prince_rounds_sub_Result_s2[30]), .ZN(prince_rounds_sub_Result_s2[28])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s2_U1 ( .A(
        prince_rounds_sub_Result_s2[29]), .B(
        prince_rounds_sub_Inv_Result_s2[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s2_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s3_U4 ( .A(
        prince_rounds_sub_Inv_Result_s3[30]), .ZN(
        prince_rounds_sub_Result_s3[31]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s3_n5), .B(
        prince_rounds_sub_Result_s3[29]), .ZN(prince_rounds_sub_Result_s3[28])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s3_U2 ( .A(
        prince_rounds_sub_Result_s3[30]), .B(
        prince_rounds_sub_Inv_Result_s3[29]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s3_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_7_A_inst_s3_U1 ( .A(
        prince_rounds_sub_Inv_Result_s3[28]), .ZN(
        prince_rounds_sub_Result_s3[29]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s1_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[35]), .B(
        prince_rounds_SR_Result_s1[18]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s1_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[32]), .B(
        prince_rounds_SR_Result_s1[17]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s1_n21), .B(
        prince_rounds_SR_Result_s1[16]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s1_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s1[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s1_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s1_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[35]), .B(
        prince_rounds_round_inputXORkeyRCON_s1[32]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s1_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[34]), .B(
        prince_rounds_SR_Result_s1[19]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_InAffin_s1_3_) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_U8 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[34]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_InAffin_s2_3_) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_U7 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[19]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[35]), .B(
        prince_rounds_SR_Result_s2[18]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2[2]) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_U5 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[32]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_U4 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_n16), .B(
        prince_rounds_SR_Result_s2[16]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[33]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_n16) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[35]), .B(
        prince_rounds_round_inputXORkeyRCON_s2[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s2_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s3_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[35]), .B(
        prince_rounds_SR_Result_s3[18]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s3_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[32]), .B(
        prince_rounds_SR_Result_s3[17]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s3_n21), .B(
        prince_rounds_SR_Result_s3[16]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s3_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s3[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s3_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s3_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[35]), .B(
        prince_rounds_round_inputXORkeyRCON_s3[32]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s3_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_Pass_inst_s3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[34]), .B(
        prince_rounds_SR_Result_s3[19]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_InAffin_s3_3_) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[3]), .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_InAffin_s1_3_), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_InAffin_s2_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_InAffin_s3_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[2]), .B(
        r[36]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_n3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[3]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3[0]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_1__CF_Inst_U1 ( 
        .A(r[0]), .B(r[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_2__CF_Inst_U1 ( 
        .A(r[1]), .B(r[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_4__CF_Inst_U1 ( 
        .A(r[2]), .B(r[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_5__CF_Inst_U1 ( 
        .A(r[3]), .B(r[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_7__CF_Inst_U1 ( 
        .A(r[4]), .B(r[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_8__CF_Inst_U1 ( 
        .A(r[5]), .B(r[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_11__CF_Inst_U1 ( 
        .A(r[7]), .B(r[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_14__CF_Inst_U1 ( 
        .A(r[9]), .B(r[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_16__CF_Inst_U1 ( 
        .A(r[10]), .B(r[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_17__CF_Inst_U1 ( 
        .A(r[11]), .B(r[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_1_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_1_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst1_InstXOR_1__Compression3_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_1_out1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1[2]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_1_out1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[2]), .B(r[37]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_2_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_2_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_2_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_1__CF_Inst_U1 ( 
        .A(r[12]), .B(r[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_2__CF_Inst_U1 ( 
        .A(r[13]), .B(r[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_4__CF_Inst_U1 ( 
        .A(r[14]), .B(r[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_5__CF_Inst_U1 ( 
        .A(r[15]), .B(r[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_7__CF_Inst_U1 ( 
        .A(r[16]), .B(r[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_8__CF_Inst_U1 ( 
        .A(r[17]), .B(r[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_10__CF_Inst_U1 ( 
        .A(r[18]), .B(r[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_11__CF_Inst_U1 ( 
        .A(r[19]), .B(r[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_13__CF_Inst_U1 ( 
        .A(r[20]), .B(r[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_14__CF_Inst_U1 ( 
        .A(r[21]), .B(r[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_16__CF_Inst_U1 ( 
        .A(r[22]), .B(r[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_17__CF_Inst_U1 ( 
        .A(r[23]), .B(r[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_2_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_2_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_2_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst2_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_2_out1[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_2_out1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2Affine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_2_out2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2Affine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_2_out2[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2Affine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_2_out3[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2Affine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_2_out3[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[2]), .B(1'b0), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s1[34]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s2[34]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s3[34]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_1__CF_Inst_U1 ( 
        .A(r[24]), .B(r[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_2__CF_Inst_U1 ( 
        .A(r[25]), .B(r[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_4__CF_Inst_U1 ( 
        .A(r[26]), .B(r[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_5__CF_Inst_U1 ( 
        .A(r[27]), .B(r[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_7__CF_Inst_U1 ( 
        .A(r[28]), .B(r[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_8__CF_Inst_U1 ( 
        .A(r[29]), .B(r[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_10__CF_Inst_U1 ( 
        .A(r[30]), .B(r[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_11__CF_Inst_U1 ( 
        .A(r[31]), .B(r[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_13__CF_Inst_U1 ( 
        .A(r[32]), .B(r[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_14__CF_Inst_U1 ( 
        .A(r[33]), .B(r[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_16__CF_Inst_U1 ( 
        .A(r[34]), .B(r[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_17__CF_Inst_U1 ( 
        .A(r[35]), .B(r[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_inst3_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_OutputAffine1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out1[3]), .Z(
        prince_rounds_sub_Result_s1[35]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_OutputAffine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out1[0]), .B(
        prince_rounds_sub_Result_s1[34]), .ZN(
        prince_rounds_sub_Inv_Result_s1[33]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_OutputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out1[0]), .Z(
        prince_rounds_sub_Result_s1[33]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_OutputAffine2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out2[3]), .Z(
        prince_rounds_sub_Result_s2[35]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_OutputAffine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out2[0]), .B(
        prince_rounds_sub_Result_s2[34]), .Z(
        prince_rounds_sub_Inv_Result_s2[33]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_OutputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out2[0]), .Z(
        prince_rounds_sub_Result_s2[33]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_OutputAffine3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out3[3]), .Z(
        prince_rounds_sub_Inv_Result_s3[34]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_OutputAffine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out3[0]), .B(
        prince_rounds_sub_Result_s3[34]), .Z(
        prince_rounds_sub_Inv_Result_s3[33]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_OutputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_8_Sub_Q294_3_out3[0]), .Z(
        prince_rounds_sub_Inv_Result_s3[32]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s1_n3), .B(
        prince_rounds_sub_Result_s1[34]), .ZN(prince_rounds_sub_Result_s1[32])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s1_U1 ( .A(
        prince_rounds_sub_Result_s1[33]), .B(
        prince_rounds_sub_Inv_Result_s1[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s2_n3), .B(
        prince_rounds_sub_Result_s2[34]), .ZN(prince_rounds_sub_Result_s2[32])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s2_U1 ( .A(
        prince_rounds_sub_Result_s2[33]), .B(
        prince_rounds_sub_Inv_Result_s2[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s2_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s3_U4 ( .A(
        prince_rounds_sub_Inv_Result_s3[34]), .ZN(
        prince_rounds_sub_Result_s3[35]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s3_n5), .B(
        prince_rounds_sub_Result_s3[33]), .ZN(prince_rounds_sub_Result_s3[32])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s3_U2 ( .A(
        prince_rounds_sub_Result_s3[34]), .B(
        prince_rounds_sub_Inv_Result_s3[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s3_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_8_A_inst_s3_U1 ( .A(
        prince_rounds_sub_Inv_Result_s3[32]), .ZN(
        prince_rounds_sub_Result_s3[33]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s1_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[39]), .B(
        prince_rounds_SR_Result_s1[6]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s1_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[36]), .B(
        prince_rounds_SR_Result_s1[5]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s1_n21), .B(
        prince_rounds_SR_Result_s1[4]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s1_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s1[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s1_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s1_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[39]), .B(
        prince_rounds_round_inputXORkeyRCON_s1[36]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s1_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[38]), .B(
        prince_rounds_SR_Result_s1[7]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_InAffin_s1_3_) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_U8 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[38]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_InAffin_s2_3_) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_U7 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[7]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[39]), .B(
        prince_rounds_SR_Result_s2[6]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2[2]) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_U5 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[36]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_U4 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_n16), .B(
        prince_rounds_SR_Result_s2[4]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[37]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_n16) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[39]), .B(
        prince_rounds_round_inputXORkeyRCON_s2[36]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s2_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s3_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[39]), .B(
        prince_rounds_SR_Result_s3[6]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s3_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[36]), .B(
        prince_rounds_SR_Result_s3[5]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s3_n19), .B(
        prince_rounds_SR_Result_s3[4]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s3_n18), .B(
        prince_rounds_round_inputXORkeyRCON_s3[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s3_n19) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s3_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[39]), .B(
        prince_rounds_round_inputXORkeyRCON_s3[36]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s3_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_Pass_inst_s3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[38]), .B(
        prince_rounds_SR_Result_s3[7]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_InAffin_s3_3_) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1[0]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1[1]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1[2]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1[3]), .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1[0]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1[1]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[1]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1[2]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[2]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1[3]), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[3]), .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_InAffin_s1_3_), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_InAffin_s2_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_InAffin_s3_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[2]), .B(
        r[36]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_n3)
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2[0]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[3]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3[0]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_1__CF_Inst_U1 ( 
        .A(r[0]), .B(r[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_2__CF_Inst_U1 ( 
        .A(r[1]), .B(r[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_4__CF_Inst_U1 ( 
        .A(r[2]), .B(r[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_5__CF_Inst_U1 ( 
        .A(r[3]), .B(r[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_7__CF_Inst_U1 ( 
        .A(r[4]), .B(r[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_8__CF_Inst_U1 ( 
        .A(r[5]), .B(r[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_11__CF_Inst_U1 ( 
        .A(r[7]), .B(r[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_14__CF_Inst_U1 ( 
        .A(r[9]), .B(r[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_16__CF_Inst_U1 ( 
        .A(r[10]), .B(r[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_17__CF_Inst_U1 ( 
        .A(r[11]), .B(r[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_1_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_1_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst1_InstXOR_1__Compression3_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_1_out1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1[2]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_1_out1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[2]), .B(r[37]), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_2_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_2_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_2_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_1__CF_Inst_U1 ( 
        .A(r[12]), .B(r[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_2__CF_Inst_U1 ( 
        .A(r[13]), .B(r[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_4__CF_Inst_U1 ( 
        .A(r[14]), .B(r[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_5__CF_Inst_U1 ( 
        .A(r[15]), .B(r[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_7__CF_Inst_U1 ( 
        .A(r[16]), .B(r[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_8__CF_Inst_U1 ( 
        .A(r[17]), .B(r[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_10__CF_Inst_U1 ( 
        .A(r[18]), .B(r[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_11__CF_Inst_U1 ( 
        .A(r[19]), .B(r[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_13__CF_Inst_U1 ( 
        .A(r[20]), .B(r[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_14__CF_Inst_U1 ( 
        .A(r[21]), .B(r[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_16__CF_Inst_U1 ( 
        .A(r[22]), .B(r[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_17__CF_Inst_U1 ( 
        .A(r[23]), .B(r[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_2_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_2_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_2_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst2_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_2_out1[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_2_out1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2Affine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_2_out2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2Affine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_2_out2[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2Affine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_2_out3[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2Affine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_2_out3[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[2]), .B(1'b0), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s1[38]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s2[38]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s3[38]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_N0), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out1[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_N1), .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out2[3]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_1__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_1__CF_Inst_U1 ( 
        .A(r[24]), .B(r[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_2__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_2__CF_Inst_U1 ( 
        .A(r[25]), .B(r[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_4__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_4__CF_Inst_U1 ( 
        .A(r[26]), .B(r[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_5__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_5__CF_Inst_U1 ( 
        .A(r[27]), .B(r[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_7__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_7__CF_Inst_U1 ( 
        .A(r[28]), .B(r[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_8__CF_Inst_n6), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_8__CF_Inst_U1 ( 
        .A(r[29]), .B(r[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_10__CF_Inst_U1 ( 
        .A(r[30]), .B(r[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_11__CF_Inst_U1 ( 
        .A(r[31]), .B(r[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_13__CF_Inst_U1 ( 
        .A(r[32]), .B(r[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_14__CF_Inst_U1 ( 
        .A(r[33]), .B(r[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_16__CF_Inst_U1 ( 
        .A(r[34]), .B(r[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_17__CF_Inst_U1 ( 
        .A(r[35]), .B(r[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_inst3_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_OutputAffine1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out1[3]), .Z(
        prince_rounds_sub_Result_s1[39]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_OutputAffine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out1[0]), .B(
        prince_rounds_sub_Result_s1[38]), .ZN(
        prince_rounds_sub_Inv_Result_s1[37]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_OutputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out1[0]), .Z(
        prince_rounds_sub_Result_s1[37]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_OutputAffine2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out2[3]), .Z(
        prince_rounds_sub_Result_s2[39]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_OutputAffine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out2[0]), .B(
        prince_rounds_sub_Result_s2[38]), .Z(
        prince_rounds_sub_Inv_Result_s2[37]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_OutputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out2[0]), .Z(
        prince_rounds_sub_Result_s2[37]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_OutputAffine3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out3[3]), .Z(
        prince_rounds_sub_Inv_Result_s3[38]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_OutputAffine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out3[0]), .B(
        prince_rounds_sub_Result_s3[38]), .Z(
        prince_rounds_sub_Inv_Result_s3[37]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_OutputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_9_Sub_Q294_3_out3[0]), .Z(
        prince_rounds_sub_Inv_Result_s3[36]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s1_n3), .B(
        prince_rounds_sub_Result_s1[38]), .ZN(prince_rounds_sub_Result_s1[36])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s1_U1 ( .A(
        prince_rounds_sub_Result_s1[37]), .B(
        prince_rounds_sub_Inv_Result_s1[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s2_n3), .B(
        prince_rounds_sub_Result_s2[38]), .ZN(prince_rounds_sub_Result_s2[36])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s2_U1 ( .A(
        prince_rounds_sub_Result_s2[37]), .B(
        prince_rounds_sub_Inv_Result_s2[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s2_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s3_U4 ( .A(
        prince_rounds_sub_Inv_Result_s3[38]), .ZN(
        prince_rounds_sub_Result_s3[39]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s3_n5), .B(
        prince_rounds_sub_Result_s3[37]), .ZN(prince_rounds_sub_Result_s3[36])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s3_U2 ( .A(
        prince_rounds_sub_Result_s3[38]), .B(
        prince_rounds_sub_Inv_Result_s3[37]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s3_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_9_A_inst_s3_U1 ( .A(
        prince_rounds_sub_Inv_Result_s3[36]), .ZN(
        prince_rounds_sub_Result_s3[37]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s1_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[43]), .B(
        prince_rounds_SR_Result_s1[58]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s1_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[40]), .B(
        prince_rounds_SR_Result_s1[57]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s1_n19), .B(
        prince_rounds_SR_Result_s1[56]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s1_n18), .B(
        prince_rounds_round_inputXORkeyRCON_s1[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s1_n19) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s1_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[43]), .B(
        prince_rounds_round_inputXORkeyRCON_s1[40]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s1_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[42]), .B(
        prince_rounds_SR_Result_s1[59]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_InAffin_s1_3_) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_U8 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[42]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_InAffin_s2_3_) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_U7 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[59]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[43]), .B(
        prince_rounds_SR_Result_s2[58]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2[2]) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_U5 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[40]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_U4 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_n16), .B(
        prince_rounds_SR_Result_s2[56]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[41]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_n16) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[43]), .B(
        prince_rounds_round_inputXORkeyRCON_s2[40]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s2_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s3_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[43]), .B(
        prince_rounds_SR_Result_s3[58]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s3_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[40]), .B(
        prince_rounds_SR_Result_s3[57]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s3_n19), .B(
        prince_rounds_SR_Result_s3[56]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s3_n18), .B(
        prince_rounds_round_inputXORkeyRCON_s3[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s3_n19) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s3_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[43]), .B(
        prince_rounds_round_inputXORkeyRCON_s3[40]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s3_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_Pass_inst_s3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[42]), .B(
        prince_rounds_SR_Result_s3[59]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_InAffin_s3_3_) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[3]), .QN()
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_InAffin_s1_3_), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_InAffin_s2_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_InAffin_s3_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[2]), .B(
        r[36]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[3]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3[0]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_1__CF_Inst_U1 ( 
        .A(r[0]), .B(r[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_2__CF_Inst_U1 ( 
        .A(r[1]), .B(r[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_4__CF_Inst_U1 ( 
        .A(r[2]), .B(r[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_5__CF_Inst_U1 ( 
        .A(r[3]), .B(r[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_7__CF_Inst_U1 ( 
        .A(r[4]), .B(r[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_8__CF_Inst_U1 ( 
        .A(r[5]), .B(r[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_11__CF_Inst_U1 ( 
        .A(r[7]), .B(r[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_14__CF_Inst_U1 ( 
        .A(r[9]), .B(r[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_16__CF_Inst_U1 ( 
        .A(r[10]), .B(r[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_17__CF_Inst_U1 ( 
        .A(r[11]), .B(r[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_1_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_1_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst1_InstXOR_1__Compression3_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_1_out1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1[2]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_1_out1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[2]), .B(r[37]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_2_out1[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_2_out2[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_2_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_1__CF_Inst_U1 ( 
        .A(r[12]), .B(r[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_2__CF_Inst_U1 ( 
        .A(r[13]), .B(r[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_4__CF_Inst_U1 ( 
        .A(r[14]), .B(r[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_5__CF_Inst_U1 ( 
        .A(r[15]), .B(r[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_7__CF_Inst_U1 ( 
        .A(r[16]), .B(r[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_8__CF_Inst_U1 ( 
        .A(r[17]), .B(r[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_10__CF_Inst_U1 ( 
        .A(r[18]), .B(r[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_11__CF_Inst_U1 ( 
        .A(r[19]), .B(r[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_13__CF_Inst_U1 ( 
        .A(r[20]), .B(r[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_14__CF_Inst_U1 ( 
        .A(r[21]), .B(r[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_16__CF_Inst_U1 ( 
        .A(r[22]), .B(r[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_17__CF_Inst_U1 ( 
        .A(r[23]), .B(r[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_2_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_2_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_2_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst2_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_2_out1[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_2_out1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2Affine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_2_out2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2Affine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_2_out2[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2Affine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_2_out3[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2Affine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_2_out3[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[2]), .B(1'b0), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s1[42]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s2[42]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s3[42]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out1[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out2[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_1__CF_Inst_U1 ( 
        .A(r[24]), .B(r[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_2__CF_Inst_U1 ( 
        .A(r[25]), .B(r[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_4__CF_Inst_U1 ( 
        .A(r[26]), .B(r[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_5__CF_Inst_U1 ( 
        .A(r[27]), .B(r[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_7__CF_Inst_U1 ( 
        .A(r[28]), .B(r[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_8__CF_Inst_U1 ( 
        .A(r[29]), .B(r[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_10__CF_Inst_U1 ( 
        .A(r[30]), .B(r[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_11__CF_Inst_U1 ( 
        .A(r[31]), .B(r[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_13__CF_Inst_U1 ( 
        .A(r[32]), .B(r[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_14__CF_Inst_U1 ( 
        .A(r[33]), .B(r[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_16__CF_Inst_U1 ( 
        .A(r[34]), .B(r[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_17__CF_Inst_U1 ( 
        .A(r[35]), .B(r[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_inst3_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_OutputAffine1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out1[3]), .Z(
        prince_rounds_sub_Result_s1[43]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_OutputAffine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out1[0]), .B(
        prince_rounds_sub_Result_s1[42]), .ZN(
        prince_rounds_sub_Inv_Result_s1[41]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_OutputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out1[0]), .Z(
        prince_rounds_sub_Result_s1[41]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_OutputAffine2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out2[3]), .Z(
        prince_rounds_sub_Result_s2[43]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_OutputAffine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out2[0]), .B(
        prince_rounds_sub_Result_s2[42]), .Z(
        prince_rounds_sub_Inv_Result_s2[41]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_OutputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out2[0]), .Z(
        prince_rounds_sub_Result_s2[41]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_OutputAffine3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out3[3]), .Z(
        prince_rounds_sub_Inv_Result_s3[42]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_OutputAffine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out3[0]), .B(
        prince_rounds_sub_Result_s3[42]), .Z(
        prince_rounds_sub_Inv_Result_s3[41]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_OutputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_10_Sub_Q294_3_out3[0]), .Z(
        prince_rounds_sub_Inv_Result_s3[40]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s1_n3), .B(
        prince_rounds_sub_Result_s1[42]), .ZN(prince_rounds_sub_Result_s1[40])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s1_U1 ( .A(
        prince_rounds_sub_Result_s1[41]), .B(
        prince_rounds_sub_Inv_Result_s1[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s2_n3), .B(
        prince_rounds_sub_Result_s2[42]), .ZN(prince_rounds_sub_Result_s2[40])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s2_U1 ( .A(
        prince_rounds_sub_Result_s2[41]), .B(
        prince_rounds_sub_Inv_Result_s2[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s2_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s3_U4 ( .A(
        prince_rounds_sub_Inv_Result_s3[42]), .ZN(
        prince_rounds_sub_Result_s3[43]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s3_n5), .B(
        prince_rounds_sub_Result_s3[41]), .ZN(prince_rounds_sub_Result_s3[40])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s3_U2 ( .A(
        prince_rounds_sub_Result_s3[42]), .B(
        prince_rounds_sub_Inv_Result_s3[41]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s3_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_10_A_inst_s3_U1 ( .A(
        prince_rounds_sub_Inv_Result_s3[40]), .ZN(
        prince_rounds_sub_Result_s3[41]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s1_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[47]), .B(
        prince_rounds_SR_Result_s1[46]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s1_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[44]), .B(
        prince_rounds_SR_Result_s1[45]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s1_n19), .B(
        prince_rounds_SR_Result_s1[44]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s1_n18), .B(
        prince_rounds_round_inputXORkeyRCON_s1[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s1_n19) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s1_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[47]), .B(
        prince_rounds_round_inputXORkeyRCON_s1[44]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s1_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[46]), .B(
        prince_rounds_SR_Result_s1[47]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_InAffin_s1_3_) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_U8 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[46]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_InAffin_s2_3_) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_U7 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[47]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[47]), .B(
        prince_rounds_SR_Result_s2[46]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2[2]) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_U5 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[44]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_U4 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_n16), .B(
        prince_rounds_SR_Result_s2[44]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[45]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_n16) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[47]), .B(
        prince_rounds_round_inputXORkeyRCON_s2[44]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s2_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s3_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[47]), .B(
        prince_rounds_SR_Result_s3[46]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s3_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[44]), .B(
        prince_rounds_SR_Result_s3[45]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s3_n19), .B(
        prince_rounds_SR_Result_s3[44]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s3_n18), .B(
        prince_rounds_round_inputXORkeyRCON_s3[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s3_n19) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s3_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[47]), .B(
        prince_rounds_round_inputXORkeyRCON_s3[44]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s3_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_Pass_inst_s3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[46]), .B(
        prince_rounds_SR_Result_s3[47]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_InAffin_s3_3_) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[3]), .QN()
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_InAffin_s1_3_), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_InAffin_s2_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_InAffin_s3_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[2]), .B(
        r[36]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[3]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3[0]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_1__CF_Inst_U1 ( 
        .A(r[0]), .B(r[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_2__CF_Inst_U1 ( 
        .A(r[1]), .B(r[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_4__CF_Inst_U1 ( 
        .A(r[2]), .B(r[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_5__CF_Inst_U1 ( 
        .A(r[3]), .B(r[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_7__CF_Inst_U1 ( 
        .A(r[4]), .B(r[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_8__CF_Inst_U1 ( 
        .A(r[5]), .B(r[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_11__CF_Inst_U1 ( 
        .A(r[7]), .B(r[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_14__CF_Inst_U1 ( 
        .A(r[9]), .B(r[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_16__CF_Inst_U1 ( 
        .A(r[10]), .B(r[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_17__CF_Inst_U1 ( 
        .A(r[11]), .B(r[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_1_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_1_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst1_InstXOR_1__Compression3_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_1_out1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1[2]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_1_out1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[2]), .B(r[37]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_2_out1[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_2_out2[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_2_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_1__CF_Inst_U1 ( 
        .A(r[12]), .B(r[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_2__CF_Inst_U1 ( 
        .A(r[13]), .B(r[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_4__CF_Inst_U1 ( 
        .A(r[14]), .B(r[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_5__CF_Inst_U1 ( 
        .A(r[15]), .B(r[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_7__CF_Inst_U1 ( 
        .A(r[16]), .B(r[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_8__CF_Inst_U1 ( 
        .A(r[17]), .B(r[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_10__CF_Inst_U1 ( 
        .A(r[18]), .B(r[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_11__CF_Inst_U1 ( 
        .A(r[19]), .B(r[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_13__CF_Inst_U1 ( 
        .A(r[20]), .B(r[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_14__CF_Inst_U1 ( 
        .A(r[21]), .B(r[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_16__CF_Inst_U1 ( 
        .A(r[22]), .B(r[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_17__CF_Inst_U1 ( 
        .A(r[23]), .B(r[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_2_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_2_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_2_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst2_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_2_out1[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_2_out1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2Affine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_2_out2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2Affine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_2_out2[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2Affine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_2_out3[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2Affine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_2_out3[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[2]), .B(1'b0), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s1[46]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s2[46]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s3[46]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out1[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out2[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_1__CF_Inst_U1 ( 
        .A(r[24]), .B(r[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_2__CF_Inst_U1 ( 
        .A(r[25]), .B(r[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_4__CF_Inst_U1 ( 
        .A(r[26]), .B(r[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_5__CF_Inst_U1 ( 
        .A(r[27]), .B(r[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_7__CF_Inst_U1 ( 
        .A(r[28]), .B(r[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_8__CF_Inst_U1 ( 
        .A(r[29]), .B(r[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_10__CF_Inst_U1 ( 
        .A(r[30]), .B(r[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_11__CF_Inst_U1 ( 
        .A(r[31]), .B(r[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_13__CF_Inst_U1 ( 
        .A(r[32]), .B(r[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_14__CF_Inst_U1 ( 
        .A(r[33]), .B(r[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_16__CF_Inst_U1 ( 
        .A(r[34]), .B(r[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_17__CF_Inst_U1 ( 
        .A(r[35]), .B(r[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_inst3_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_OutputAffine1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out1[3]), .Z(
        prince_rounds_sub_Result_s1[47]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_OutputAffine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out1[0]), .B(
        prince_rounds_sub_Result_s1[46]), .ZN(
        prince_rounds_sub_Inv_Result_s1[45]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_OutputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out1[0]), .Z(
        prince_rounds_sub_Result_s1[45]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_OutputAffine2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out2[3]), .Z(
        prince_rounds_sub_Result_s2[47]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_OutputAffine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out2[0]), .B(
        prince_rounds_sub_Result_s2[46]), .Z(
        prince_rounds_sub_Inv_Result_s2[45]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_OutputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out2[0]), .Z(
        prince_rounds_sub_Result_s2[45]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_OutputAffine3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out3[3]), .Z(
        prince_rounds_sub_Inv_Result_s3[46]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_OutputAffine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out3[0]), .B(
        prince_rounds_sub_Result_s3[46]), .Z(
        prince_rounds_sub_Inv_Result_s3[45]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_OutputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_11_Sub_Q294_3_out3[0]), .Z(
        prince_rounds_sub_Inv_Result_s3[44]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s1_n3), .B(
        prince_rounds_sub_Result_s1[46]), .ZN(prince_rounds_sub_Result_s1[44])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s1_U1 ( .A(
        prince_rounds_sub_Result_s1[45]), .B(
        prince_rounds_sub_Inv_Result_s1[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s2_n3), .B(
        prince_rounds_sub_Result_s2[46]), .ZN(prince_rounds_sub_Result_s2[44])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s2_U1 ( .A(
        prince_rounds_sub_Result_s2[45]), .B(
        prince_rounds_sub_Inv_Result_s2[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s2_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s3_U4 ( .A(
        prince_rounds_sub_Inv_Result_s3[46]), .ZN(
        prince_rounds_sub_Result_s3[47]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s3_n5), .B(
        prince_rounds_sub_Result_s3[45]), .ZN(prince_rounds_sub_Result_s3[44])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s3_U2 ( .A(
        prince_rounds_sub_Result_s3[46]), .B(
        prince_rounds_sub_Inv_Result_s3[45]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s3_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_11_A_inst_s3_U1 ( .A(
        prince_rounds_sub_Inv_Result_s3[44]), .ZN(
        prince_rounds_sub_Result_s3[45]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s1_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[51]), .B(
        prince_rounds_SR_Result_s1[34]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s1_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[48]), .B(
        prince_rounds_SR_Result_s1[33]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s1_n19), .B(
        prince_rounds_SR_Result_s1[32]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s1_n18), .B(
        prince_rounds_round_inputXORkeyRCON_s1[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s1_n19) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s1_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[51]), .B(
        prince_rounds_round_inputXORkeyRCON_s1[48]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s1_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[50]), .B(
        prince_rounds_SR_Result_s1[35]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_InAffin_s1_3_) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_U8 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[50]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_InAffin_s2_3_) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_U7 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[35]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[51]), .B(
        prince_rounds_SR_Result_s2[34]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2[2]) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_U5 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[48]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_U4 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[33]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_n16), .B(
        prince_rounds_SR_Result_s2[32]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[49]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_n16) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[51]), .B(
        prince_rounds_round_inputXORkeyRCON_s2[48]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s2_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s3_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[51]), .B(
        prince_rounds_SR_Result_s3[34]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s3_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[48]), .B(
        prince_rounds_SR_Result_s3[33]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s3_n19), .B(
        prince_rounds_SR_Result_s3[32]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s3_n18), .B(
        prince_rounds_round_inputXORkeyRCON_s3[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s3_n19) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s3_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[51]), .B(
        prince_rounds_round_inputXORkeyRCON_s3[48]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s3_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_Pass_inst_s3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[50]), .B(
        prince_rounds_SR_Result_s3[35]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_InAffin_s3_3_) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[3]), .QN()
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_InAffin_s1_3_), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_InAffin_s2_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_InAffin_s3_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[2]), .B(
        r[36]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[3]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3[0]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_1__CF_Inst_U1 ( 
        .A(r[0]), .B(r[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_2__CF_Inst_U1 ( 
        .A(r[1]), .B(r[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_4__CF_Inst_U1 ( 
        .A(r[2]), .B(r[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_5__CF_Inst_U1 ( 
        .A(r[3]), .B(r[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_7__CF_Inst_U1 ( 
        .A(r[4]), .B(r[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_8__CF_Inst_U1 ( 
        .A(r[5]), .B(r[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_11__CF_Inst_U1 ( 
        .A(r[7]), .B(r[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_14__CF_Inst_U1 ( 
        .A(r[9]), .B(r[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_16__CF_Inst_U1 ( 
        .A(r[10]), .B(r[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_17__CF_Inst_U1 ( 
        .A(r[11]), .B(r[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_1_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_1_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst1_InstXOR_1__Compression3_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_1_out1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1[2]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_1_out1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[2]), .B(r[37]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_2_out1[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_2_out2[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_2_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_1__CF_Inst_U1 ( 
        .A(r[12]), .B(r[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_2__CF_Inst_U1 ( 
        .A(r[13]), .B(r[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_4__CF_Inst_U1 ( 
        .A(r[14]), .B(r[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_5__CF_Inst_U1 ( 
        .A(r[15]), .B(r[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_7__CF_Inst_U1 ( 
        .A(r[16]), .B(r[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_8__CF_Inst_U1 ( 
        .A(r[17]), .B(r[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_10__CF_Inst_U1 ( 
        .A(r[18]), .B(r[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_11__CF_Inst_U1 ( 
        .A(r[19]), .B(r[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_13__CF_Inst_U1 ( 
        .A(r[20]), .B(r[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_14__CF_Inst_U1 ( 
        .A(r[21]), .B(r[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_16__CF_Inst_U1 ( 
        .A(r[22]), .B(r[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_17__CF_Inst_U1 ( 
        .A(r[23]), .B(r[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_2_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_2_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_2_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst2_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_2_out1[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_2_out1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2Affine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_2_out2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2Affine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_2_out2[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2Affine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_2_out3[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2Affine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_2_out3[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[2]), .B(1'b0), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s1[50]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s2[50]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s3[50]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out1[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out2[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_1__CF_Inst_U1 ( 
        .A(r[24]), .B(r[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_2__CF_Inst_U1 ( 
        .A(r[25]), .B(r[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_4__CF_Inst_U1 ( 
        .A(r[26]), .B(r[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_5__CF_Inst_U1 ( 
        .A(r[27]), .B(r[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_7__CF_Inst_U1 ( 
        .A(r[28]), .B(r[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_8__CF_Inst_U1 ( 
        .A(r[29]), .B(r[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_10__CF_Inst_U1 ( 
        .A(r[30]), .B(r[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_11__CF_Inst_U1 ( 
        .A(r[31]), .B(r[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_13__CF_Inst_U1 ( 
        .A(r[32]), .B(r[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_14__CF_Inst_U1 ( 
        .A(r[33]), .B(r[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_16__CF_Inst_U1 ( 
        .A(r[34]), .B(r[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_17__CF_Inst_U1 ( 
        .A(r[35]), .B(r[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_inst3_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_OutputAffine1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out1[3]), .Z(
        prince_rounds_sub_Result_s1[51]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_OutputAffine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out1[0]), .B(
        prince_rounds_sub_Result_s1[50]), .ZN(
        prince_rounds_sub_Inv_Result_s1[49]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_OutputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out1[0]), .Z(
        prince_rounds_sub_Result_s1[49]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_OutputAffine2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out2[3]), .Z(
        prince_rounds_sub_Result_s2[51]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_OutputAffine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out2[0]), .B(
        prince_rounds_sub_Result_s2[50]), .Z(
        prince_rounds_sub_Inv_Result_s2[49]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_OutputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out2[0]), .Z(
        prince_rounds_sub_Result_s2[49]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_OutputAffine3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out3[3]), .Z(
        prince_rounds_sub_Inv_Result_s3[50]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_OutputAffine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out3[0]), .B(
        prince_rounds_sub_Result_s3[50]), .Z(
        prince_rounds_sub_Inv_Result_s3[49]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_OutputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_12_Sub_Q294_3_out3[0]), .Z(
        prince_rounds_sub_Inv_Result_s3[48]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s1_n3), .B(
        prince_rounds_sub_Result_s1[50]), .ZN(prince_rounds_sub_Result_s1[48])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s1_U1 ( .A(
        prince_rounds_sub_Result_s1[49]), .B(
        prince_rounds_sub_Inv_Result_s1[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s2_n3), .B(
        prince_rounds_sub_Result_s2[50]), .ZN(prince_rounds_sub_Result_s2[48])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s2_U1 ( .A(
        prince_rounds_sub_Result_s2[49]), .B(
        prince_rounds_sub_Inv_Result_s2[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s2_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s3_U4 ( .A(
        prince_rounds_sub_Inv_Result_s3[50]), .ZN(
        prince_rounds_sub_Result_s3[51]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s3_n5), .B(
        prince_rounds_sub_Result_s3[49]), .ZN(prince_rounds_sub_Result_s3[48])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s3_U2 ( .A(
        prince_rounds_sub_Result_s3[50]), .B(
        prince_rounds_sub_Inv_Result_s3[49]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s3_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_12_A_inst_s3_U1 ( .A(
        prince_rounds_sub_Inv_Result_s3[48]), .ZN(
        prince_rounds_sub_Result_s3[49]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s1_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[55]), .B(
        prince_rounds_SR_Result_s1[22]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s1_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[52]), .B(
        prince_rounds_SR_Result_s1[21]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s1_n21), .B(
        prince_rounds_SR_Result_s1[20]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s1_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s1[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s1_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s1_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[55]), .B(
        prince_rounds_round_inputXORkeyRCON_s1[52]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s1_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[54]), .B(
        prince_rounds_SR_Result_s1[23]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_InAffin_s1_3_) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_U8 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[54]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_InAffin_s2_3_) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_U7 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[23]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[55]), .B(
        prince_rounds_SR_Result_s2[22]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2[2]) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_U5 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[52]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_U4 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[21]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_n16), .B(
        prince_rounds_SR_Result_s2[20]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[53]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_n16) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[55]), .B(
        prince_rounds_round_inputXORkeyRCON_s2[52]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s2_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s3_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[55]), .B(
        prince_rounds_SR_Result_s3[22]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s3_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[52]), .B(
        prince_rounds_SR_Result_s3[21]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s3_n21), .B(
        prince_rounds_SR_Result_s3[20]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s3_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s3[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s3_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s3_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[55]), .B(
        prince_rounds_round_inputXORkeyRCON_s3[52]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s3_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_Pass_inst_s3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[54]), .B(
        prince_rounds_SR_Result_s3[23]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_InAffin_s3_3_) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[3]), .QN()
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_InAffin_s1_3_), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_InAffin_s2_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_InAffin_s3_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[2]), .B(
        r[36]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[3]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3[0]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_1__CF_Inst_U1 ( 
        .A(r[0]), .B(r[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_2__CF_Inst_U1 ( 
        .A(r[1]), .B(r[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_4__CF_Inst_U1 ( 
        .A(r[2]), .B(r[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_5__CF_Inst_U1 ( 
        .A(r[3]), .B(r[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_7__CF_Inst_U1 ( 
        .A(r[4]), .B(r[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_8__CF_Inst_U1 ( 
        .A(r[5]), .B(r[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_11__CF_Inst_U1 ( 
        .A(r[7]), .B(r[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_14__CF_Inst_U1 ( 
        .A(r[9]), .B(r[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_16__CF_Inst_U1 ( 
        .A(r[10]), .B(r[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_17__CF_Inst_U1 ( 
        .A(r[11]), .B(r[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_1_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_1_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst1_InstXOR_1__Compression3_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_1_out1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1[2]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_1_out1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[2]), .B(r[37]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_2_out1[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_2_out2[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_2_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_1__CF_Inst_U1 ( 
        .A(r[12]), .B(r[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_2__CF_Inst_U1 ( 
        .A(r[13]), .B(r[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_4__CF_Inst_U1 ( 
        .A(r[14]), .B(r[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_5__CF_Inst_U1 ( 
        .A(r[15]), .B(r[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_7__CF_Inst_U1 ( 
        .A(r[16]), .B(r[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_8__CF_Inst_U1 ( 
        .A(r[17]), .B(r[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_10__CF_Inst_U1 ( 
        .A(r[18]), .B(r[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_11__CF_Inst_U1 ( 
        .A(r[19]), .B(r[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_13__CF_Inst_U1 ( 
        .A(r[20]), .B(r[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_14__CF_Inst_U1 ( 
        .A(r[21]), .B(r[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_16__CF_Inst_U1 ( 
        .A(r[22]), .B(r[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_17__CF_Inst_U1 ( 
        .A(r[23]), .B(r[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_2_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_2_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_2_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst2_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_2_out1[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_2_out1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2Affine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_2_out2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2Affine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_2_out2[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2Affine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_2_out3[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2Affine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_2_out3[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[2]), .B(1'b0), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s1[54]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s2[54]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s3[54]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out1[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out2[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_1__CF_Inst_U1 ( 
        .A(r[24]), .B(r[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_2__CF_Inst_U1 ( 
        .A(r[25]), .B(r[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_4__CF_Inst_U1 ( 
        .A(r[26]), .B(r[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_5__CF_Inst_U1 ( 
        .A(r[27]), .B(r[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_7__CF_Inst_U1 ( 
        .A(r[28]), .B(r[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_8__CF_Inst_U1 ( 
        .A(r[29]), .B(r[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_10__CF_Inst_U1 ( 
        .A(r[30]), .B(r[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_11__CF_Inst_U1 ( 
        .A(r[31]), .B(r[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_13__CF_Inst_U1 ( 
        .A(r[32]), .B(r[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_14__CF_Inst_U1 ( 
        .A(r[33]), .B(r[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_16__CF_Inst_U1 ( 
        .A(r[34]), .B(r[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_17__CF_Inst_U1 ( 
        .A(r[35]), .B(r[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_inst3_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_OutputAffine1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out1[3]), .Z(
        prince_rounds_sub_Result_s1[55]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_OutputAffine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out1[0]), .B(
        prince_rounds_sub_Result_s1[54]), .ZN(
        prince_rounds_sub_Inv_Result_s1[53]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_OutputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out1[0]), .Z(
        prince_rounds_sub_Result_s1[53]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_OutputAffine2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out2[3]), .Z(
        prince_rounds_sub_Result_s2[55]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_OutputAffine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out2[0]), .B(
        prince_rounds_sub_Result_s2[54]), .Z(
        prince_rounds_sub_Inv_Result_s2[53]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_OutputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out2[0]), .Z(
        prince_rounds_sub_Result_s2[53]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_OutputAffine3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out3[3]), .Z(
        prince_rounds_sub_Inv_Result_s3[54]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_OutputAffine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out3[0]), .B(
        prince_rounds_sub_Result_s3[54]), .Z(
        prince_rounds_sub_Inv_Result_s3[53]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_OutputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_13_Sub_Q294_3_out3[0]), .Z(
        prince_rounds_sub_Inv_Result_s3[52]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s1_n3), .B(
        prince_rounds_sub_Result_s1[54]), .ZN(prince_rounds_sub_Result_s1[52])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s1_U1 ( .A(
        prince_rounds_sub_Result_s1[53]), .B(
        prince_rounds_sub_Inv_Result_s1[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s2_n3), .B(
        prince_rounds_sub_Result_s2[54]), .ZN(prince_rounds_sub_Result_s2[52])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s2_U1 ( .A(
        prince_rounds_sub_Result_s2[53]), .B(
        prince_rounds_sub_Inv_Result_s2[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s2_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s3_U4 ( .A(
        prince_rounds_sub_Inv_Result_s3[54]), .ZN(
        prince_rounds_sub_Result_s3[55]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s3_n5), .B(
        prince_rounds_sub_Result_s3[53]), .ZN(prince_rounds_sub_Result_s3[52])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s3_U2 ( .A(
        prince_rounds_sub_Result_s3[54]), .B(
        prince_rounds_sub_Inv_Result_s3[53]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s3_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_13_A_inst_s3_U1 ( .A(
        prince_rounds_sub_Inv_Result_s3[52]), .ZN(
        prince_rounds_sub_Result_s3[53]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s1_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[59]), .B(
        prince_rounds_SR_Result_s1[10]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s1_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[56]), .B(
        prince_rounds_SR_Result_s1[9]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s1_n21), .B(
        prince_rounds_SR_Result_s1[8]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s1_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s1[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s1_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s1_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[59]), .B(
        prince_rounds_round_inputXORkeyRCON_s1[56]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s1_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[58]), .B(
        prince_rounds_SR_Result_s1[11]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_InAffin_s1_3_) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_U8 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[58]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_InAffin_s2_3_) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_U7 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[59]), .B(
        prince_rounds_SR_Result_s2[10]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2[2]) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_U5 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[56]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_U4 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[9]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_n16), .B(
        prince_rounds_SR_Result_s2[8]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[57]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_n16) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[59]), .B(
        prince_rounds_round_inputXORkeyRCON_s2[56]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s2_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s3_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[59]), .B(
        prince_rounds_SR_Result_s3[10]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s3_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[56]), .B(
        prince_rounds_SR_Result_s3[9]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s3_n21), .B(
        prince_rounds_SR_Result_s3[8]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s3_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s3[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s3_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s3_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[59]), .B(
        prince_rounds_round_inputXORkeyRCON_s3[56]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s3_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_Pass_inst_s3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[58]), .B(
        prince_rounds_SR_Result_s3[11]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_InAffin_s3_3_) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[3]), .QN()
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_InAffin_s1_3_), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_InAffin_s2_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_InAffin_s3_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[2]), .B(
        r[36]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[3]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3[0]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_1__CF_Inst_U1 ( 
        .A(r[0]), .B(r[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_2__CF_Inst_U1 ( 
        .A(r[1]), .B(r[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_4__CF_Inst_U1 ( 
        .A(r[2]), .B(r[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_5__CF_Inst_U1 ( 
        .A(r[3]), .B(r[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_7__CF_Inst_U1 ( 
        .A(r[4]), .B(r[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_8__CF_Inst_U1 ( 
        .A(r[5]), .B(r[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_11__CF_Inst_U1 ( 
        .A(r[7]), .B(r[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_14__CF_Inst_U1 ( 
        .A(r[9]), .B(r[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_16__CF_Inst_U1 ( 
        .A(r[10]), .B(r[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_17__CF_Inst_U1 ( 
        .A(r[11]), .B(r[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_1_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_1_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst1_InstXOR_1__Compression3_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_1_out1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1[2]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_1_out1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[2]), .B(r[37]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_2_out1[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_2_out2[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_2_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_1__CF_Inst_U1 ( 
        .A(r[12]), .B(r[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_2__CF_Inst_U1 ( 
        .A(r[13]), .B(r[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_4__CF_Inst_U1 ( 
        .A(r[14]), .B(r[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_5__CF_Inst_U1 ( 
        .A(r[15]), .B(r[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_7__CF_Inst_U1 ( 
        .A(r[16]), .B(r[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_8__CF_Inst_U1 ( 
        .A(r[17]), .B(r[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_10__CF_Inst_U1 ( 
        .A(r[18]), .B(r[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_11__CF_Inst_U1 ( 
        .A(r[19]), .B(r[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_13__CF_Inst_U1 ( 
        .A(r[20]), .B(r[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_14__CF_Inst_U1 ( 
        .A(r[21]), .B(r[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_16__CF_Inst_U1 ( 
        .A(r[22]), .B(r[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_17__CF_Inst_U1 ( 
        .A(r[23]), .B(r[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_2_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_2_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_2_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst2_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_2_out1[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_2_out1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2Affine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_2_out2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2Affine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_2_out2[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2Affine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_2_out3[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2Affine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_2_out3[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[2]), .B(1'b0), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s1[58]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s2[58]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s3[58]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out1[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out2[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_1__CF_Inst_U1 ( 
        .A(r[24]), .B(r[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_2__CF_Inst_U1 ( 
        .A(r[25]), .B(r[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_4__CF_Inst_U1 ( 
        .A(r[26]), .B(r[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_5__CF_Inst_U1 ( 
        .A(r[27]), .B(r[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_7__CF_Inst_U1 ( 
        .A(r[28]), .B(r[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_8__CF_Inst_U1 ( 
        .A(r[29]), .B(r[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_10__CF_Inst_U1 ( 
        .A(r[30]), .B(r[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_11__CF_Inst_U1 ( 
        .A(r[31]), .B(r[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_13__CF_Inst_U1 ( 
        .A(r[32]), .B(r[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_14__CF_Inst_U1 ( 
        .A(r[33]), .B(r[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_16__CF_Inst_U1 ( 
        .A(r[34]), .B(r[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_17__CF_Inst_U1 ( 
        .A(r[35]), .B(r[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_inst3_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_OutputAffine1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out1[3]), .Z(
        prince_rounds_sub_Result_s1[59]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_OutputAffine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out1[0]), .B(
        prince_rounds_sub_Result_s1[58]), .ZN(
        prince_rounds_sub_Inv_Result_s1[57]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_OutputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out1[0]), .Z(
        prince_rounds_sub_Result_s1[57]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_OutputAffine2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out2[3]), .Z(
        prince_rounds_sub_Result_s2[59]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_OutputAffine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out2[0]), .B(
        prince_rounds_sub_Result_s2[58]), .Z(
        prince_rounds_sub_Inv_Result_s2[57]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_OutputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out2[0]), .Z(
        prince_rounds_sub_Result_s2[57]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_OutputAffine3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out3[3]), .Z(
        prince_rounds_sub_Inv_Result_s3[58]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_OutputAffine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out3[0]), .B(
        prince_rounds_sub_Result_s3[58]), .Z(
        prince_rounds_sub_Inv_Result_s3[57]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_OutputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_14_Sub_Q294_3_out3[0]), .Z(
        prince_rounds_sub_Inv_Result_s3[56]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s1_n3), .B(
        prince_rounds_sub_Result_s1[58]), .ZN(prince_rounds_sub_Result_s1[56])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s1_U1 ( .A(
        prince_rounds_sub_Result_s1[57]), .B(
        prince_rounds_sub_Inv_Result_s1[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s2_n3), .B(
        prince_rounds_sub_Result_s2[58]), .ZN(prince_rounds_sub_Result_s2[56])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s2_U1 ( .A(
        prince_rounds_sub_Result_s2[57]), .B(
        prince_rounds_sub_Inv_Result_s2[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s2_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s3_U4 ( .A(
        prince_rounds_sub_Inv_Result_s3[58]), .ZN(
        prince_rounds_sub_Result_s3[59]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s3_n5), .B(
        prince_rounds_sub_Result_s3[57]), .ZN(prince_rounds_sub_Result_s3[56])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s3_U2 ( .A(
        prince_rounds_sub_Result_s3[58]), .B(
        prince_rounds_sub_Inv_Result_s3[57]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s3_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_14_A_inst_s3_U1 ( .A(
        prince_rounds_sub_Inv_Result_s3[56]), .ZN(
        prince_rounds_sub_Result_s3[57]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s1_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[63]), .B(
        prince_rounds_SR_Result_s1[62]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s1_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[60]), .B(
        prince_rounds_SR_Result_s1[61]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s1_n21), .B(
        prince_rounds_SR_Result_s1[60]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s1_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s1[61]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s1_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s1_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[63]), .B(
        prince_rounds_round_inputXORkeyRCON_s1[60]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s1_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s1_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s1[62]), .B(
        prince_rounds_SR_Result_s1[63]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_InAffin_s1_3_) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_U8 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[62]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_n18), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_InAffin_s2_3_) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_U7 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[63]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_n18) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[63]), .B(
        prince_rounds_SR_Result_s2[62]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2[2]) );
  OAI21_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_U5 ( .B1(
        prince_rounds_sub_n3), .B2(prince_rounds_round_inputXORkeyRCON_s2[60]), 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_n17), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_U4 ( .A1(
        prince_rounds_sub_n3), .A2(prince_rounds_SR_Result_s2[61]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_n17) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_n16), .B(
        prince_rounds_SR_Result_s2[60]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[61]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_n15), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_n16) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s2[63]), .B(
        prince_rounds_round_inputXORkeyRCON_s2[60]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s2_n15) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s3_U6 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[63]), .B(
        prince_rounds_SR_Result_s3[62]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3[2]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s3_U5 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[60]), .B(
        prince_rounds_SR_Result_s3[61]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3[0]) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s3_n21), .B(
        prince_rounds_SR_Result_s3[60]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s3_n20), .B(
        prince_rounds_round_inputXORkeyRCON_s3[61]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s3_n21) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s3_U2 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[63]), .B(
        prince_rounds_round_inputXORkeyRCON_s3[60]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s3_n20) );
  MUX2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_Pass_inst_s3_U1 ( .A(
        prince_rounds_round_inputXORkeyRCON_s3[62]), .B(
        prince_rounds_SR_Result_s3[63]), .S(prince_rounds_sub_n3), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_InAffin_s3_3_) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg_reg_0_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1[0]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg_reg_1_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1[1]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg_reg_2_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1[2]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg_reg_3_ ( .D(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1[3]), .CK(clk), 
        .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[3]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1[0]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[0]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1[1]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[1]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1[2]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[2]), .QN()
         );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1[3]), .CK(
        clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[3]), .QN()
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_InAffin_s1_3_), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_InAffin_s2_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_InAffin_s3_3_), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[2]), .B(
        r[36]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[2]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[3]), 
        .CK(clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3[0]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_1__CF_Inst_U1 ( 
        .A(r[0]), .B(r[1]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_2__CF_Inst_U1 ( 
        .A(r[1]), .B(r[2]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_4__CF_Inst_U1 ( 
        .A(r[2]), .B(r[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_5__CF_Inst_U1 ( 
        .A(r[3]), .B(r[4]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_7__CF_Inst_U1 ( 
        .A(r[4]), .B(r[5]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[1]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_8__CF_Inst_U1 ( 
        .A(r[5]), .B(r[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_10__CF_Inst_U1 ( 
        .A(r[6]), .B(r[7]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_11__CF_Inst_U1 ( 
        .A(r[7]), .B(r[8]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_13__CF_Inst_U1 ( 
        .A(r[8]), .B(r[9]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out3_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_14__CF_Inst_U1 ( 
        .A(r[9]), .B(r[10]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_16__CF_Inst_U1 ( 
        .A(r[10]), .B(r[11]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out2_reg[2]), 
        .A2(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_InAff_out1_reg[3]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_17__CF_Inst_U1 ( 
        .A(r[11]), .B(r[6]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_1_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_1_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst1_InstXOR_1__Compression3_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_1_out1[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1[2]) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_1_out1[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1[3]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[2]), .B(r[37]), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_2_out1[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_2_out2[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_2_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_1__CF_Inst_U1 ( 
        .A(r[12]), .B(r[13]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_2__CF_Inst_U1 ( 
        .A(r[13]), .B(r[14]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_4__CF_Inst_U1 ( 
        .A(r[14]), .B(r[15]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_5__CF_Inst_U1 ( 
        .A(r[15]), .B(r[16]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_7__CF_Inst_U1 ( 
        .A(r[16]), .B(r[17]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_8__CF_Inst_U1 ( 
        .A(r[17]), .B(r[12]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_10__CF_Inst_U1 ( 
        .A(r[18]), .B(r[19]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_11__CF_Inst_U1 ( 
        .A(r[19]), .B(r[20]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_13__CF_Inst_U1 ( 
        .A(r[20]), .B(r[21]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_14__CF_Inst_U1 ( 
        .A(r[21]), .B(r[22]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_16__CF_Inst_U1 ( 
        .A(r[22]), .B(r[23]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M1_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_17__CF_Inst_U1 ( 
        .A(r[23]), .B(r[18]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_2_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_2_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_2_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3[2]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst2_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2Affine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_2_out1[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2Affine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_2_out1[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2Affine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_2_out2[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2Affine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_2_out2[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2[1]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2Affine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3[2]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_2_out3[0]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3[3]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2Affine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3[0]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_2_out3[3]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_U5 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_N1) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_U4 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[3]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_n3), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_N0) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[2]), .B(1'b0), 
        .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_n3) );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_0_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[0]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[0]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[1]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[1]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[2]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[2]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[3]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_4_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[4]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[4]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_5_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[5]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[5]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_6_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[6]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[6]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_7_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[7]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[7]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_8_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[8]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[8]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_9_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[9]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[9]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_10_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[10]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[10]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_11_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[11]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[11]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_12_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[12]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[12]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_13_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[13]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[13]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_14_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[14]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[14]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_15_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[15]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[15]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_16_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[16]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[16]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg_reg_17_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[17]), 
        .CK(clk), .Q(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[17]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_creg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s1[62]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_creg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s2[62]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_creg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[2]), .CK(
        clk), .Q(prince_rounds_sub_Result_s3[62]), .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_dreg_reg_1_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_N0), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out1[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_dreg_reg_2_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_N1), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out2[3]), 
        .QN() );
  DFF_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_dreg_reg_3_ ( 
        .D(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[3]), .CK(
        clk), .Q(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out3[3]), 
        .QN() );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_0__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_0__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[0]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_0__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_0__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_1__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_1__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_1__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[1]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_1__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_1__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_1__CF_Inst_U1 ( 
        .A(r[24]), .B(r[25]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_1__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_2__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_2__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_2__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[2]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_2__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_2__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_2__CF_Inst_U1 ( 
        .A(r[25]), .B(r[26]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_2__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_3__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_3__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[3]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_3__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_3__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_4__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_4__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_4__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[4]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_4__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_4__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_4__CF_Inst_U1 ( 
        .A(r[26]), .B(r[27]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_4__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_5__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_5__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_5__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[5]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_5__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_5__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_5__CF_Inst_U1 ( 
        .A(r[27]), .B(r[28]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_5__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_6__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_6__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[0]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[6]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_6__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_6__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_7__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_7__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_7__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[7]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_7__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_7__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_7__CF_Inst_U1 ( 
        .A(r[28]), .B(r[29]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_7__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_8__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_8__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_8__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[8]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_8__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[1]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_8__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_8__CF_Inst_U1 ( 
        .A(r[29]), .B(r[24]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_8__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_9__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_9__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[9]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_9__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_9__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_10__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_10__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_10__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[10]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_10__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_10__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_10__CF_Inst_U1 ( 
        .A(r[30]), .B(r[31]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_10__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_11__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_11__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_11__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[11]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_11__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_11__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_11__CF_Inst_U1 ( 
        .A(r[31]), .B(r[32]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_11__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_12__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_12__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[12]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_12__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_12__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_13__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_13__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_13__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[13]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_13__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_13__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_13__CF_Inst_U1 ( 
        .A(r[32]), .B(r[33]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_13__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_14__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_14__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_14__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[14]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_14__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out3_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_14__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_14__CF_Inst_U1 ( 
        .A(r[33]), .B(r[34]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_14__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_15__CF_Inst_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_15__CF_Inst_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[1]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[15]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_15__CF_Inst_U1 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_15__CF_Inst_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_16__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_16__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_16__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[16]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_16__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_16__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_16__CF_Inst_U1 ( 
        .A(r[34]), .B(r[35]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_16__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_17__CF_Inst_U3 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_17__CF_Inst_n6), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_17__CF_Inst_n5), .ZN(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Out[17]) );
  NAND2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_17__CF_Inst_U2 ( 
        .A1(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out2_reg[2]), .A2(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_M2_out1_reg[3]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_17__CF_Inst_n5) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_17__CF_Inst_U1 ( 
        .A(r[35]), .B(r[30]), .Z(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_Inst_17__CF_Inst_n6) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_0__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_0__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[2]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out1[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_0__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[0]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[1]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_0__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_0__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_0__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[5]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out2[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_0__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[3]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[4]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_0__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_0__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_0__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[8]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out3[0]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_0__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[6]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[7]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_0__Compression3_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_1__Compression1_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_1__Compression1_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[11]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out1[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_1__Compression1_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[9]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[10]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_1__Compression1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_1__Compression2_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_1__Compression2_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[14]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out2[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_1__Compression2_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[12]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[13]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_1__Compression2_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_1__Compression3_U2 ( 
        .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_1__Compression3_n3), .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[17]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out3[1]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_1__Compression3_U1 ( 
        .A(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[15]), 
        .B(prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_CF_Reg[16]), 
        .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_inst3_InstXOR_1__Compression3_n3) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_OutputAffine1_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out1[3]), .Z(
        prince_rounds_sub_Result_s1[63]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_OutputAffine1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out1[0]), .B(
        prince_rounds_sub_Result_s1[62]), .ZN(
        prince_rounds_sub_Inv_Result_s1[61]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_OutputAffine1_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out1[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out1[0]), .Z(
        prince_rounds_sub_Result_s1[61]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_OutputAffine2_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out2[3]), .Z(
        prince_rounds_sub_Result_s2[63]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_OutputAffine2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out2[0]), .B(
        prince_rounds_sub_Result_s2[62]), .Z(
        prince_rounds_sub_Inv_Result_s2[61]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_OutputAffine2_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out2[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out2[0]), .Z(
        prince_rounds_sub_Result_s2[61]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_OutputAffine3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out3[3]), .Z(
        prince_rounds_sub_Inv_Result_s3[62]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_OutputAffine3_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out3[0]), .B(
        prince_rounds_sub_Result_s3[62]), .Z(
        prince_rounds_sub_Inv_Result_s3[61]) );
  XOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_OutputAffine3_U1 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out3[1]), .B(
        prince_rounds_sub_sBoxCombined_PRINCE_15_Sub_Q294_3_out3[0]), .Z(
        prince_rounds_sub_Inv_Result_s3[60]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s1_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s1_n3), .B(
        prince_rounds_sub_Result_s1[62]), .ZN(prince_rounds_sub_Result_s1[60])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s1_U1 ( .A(
        prince_rounds_sub_Result_s1[61]), .B(
        prince_rounds_sub_Inv_Result_s1[61]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s1_n3) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s2_U2 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s2_n3), .B(
        prince_rounds_sub_Result_s2[62]), .ZN(prince_rounds_sub_Result_s2[60])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s2_U1 ( .A(
        prince_rounds_sub_Result_s2[61]), .B(
        prince_rounds_sub_Inv_Result_s2[61]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s2_n3) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s3_U4 ( .A(
        prince_rounds_sub_Inv_Result_s3[62]), .ZN(
        prince_rounds_sub_Result_s3[63]) );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s3_U3 ( .A(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s3_n5), .B(
        prince_rounds_sub_Result_s3[61]), .ZN(prince_rounds_sub_Result_s3[60])
         );
  XNOR2_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s3_U2 ( .A(
        prince_rounds_sub_Result_s3[62]), .B(
        prince_rounds_sub_Inv_Result_s3[61]), .ZN(
        prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s3_n5) );
  INV_X1 prince_rounds_sub_sBoxCombined_PRINCE_15_A_inst_s3_U1 ( .A(
        prince_rounds_sub_Inv_Result_s3[60]), .ZN(
        prince_rounds_sub_Result_s3[61]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_0_0_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_0_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_0_), .ZN(
        prince_rounds_SR_Inv_Result_s1[16]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_0_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[1]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_0_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_0_1_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_0_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_1_), .ZN(
        prince_rounds_SR_Inv_Result_s1[17]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_0_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s1[1]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_0_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_0_2_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_0_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_2_), .ZN(
        prince_rounds_SR_Inv_Result_s1[18]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_0_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[3]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_0_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_0_3_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_0_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_3_), .ZN(
        prince_rounds_SR_Inv_Result_s1[19]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_0_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[2]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_0_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_1_0_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_1_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_4_), .ZN(
        prince_rounds_SR_Inv_Result_s1[36]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_1_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[5]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_1_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_1_1_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_1_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_5_), .ZN(
        prince_rounds_SR_Inv_Result_s1[37]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_1_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s1[5]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_1_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_1_2_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_1_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_6_), .ZN(
        prince_rounds_SR_Inv_Result_s1[38]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_1_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[7]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_1_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_1_3_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_1_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_7_), .ZN(
        prince_rounds_SR_Inv_Result_s1[39]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_1_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[6]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_1_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_2_0_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_2_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_8_), .ZN(
        prince_rounds_SR_Inv_Result_s1[56]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_2_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[9]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_2_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_2_1_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_2_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_9_), .ZN(
        prince_rounds_SR_Inv_Result_s1[57]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_2_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s1[9]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_2_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_2_2_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_2_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_10_), .ZN(
        prince_rounds_SR_Inv_Result_s1[58]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_2_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[11]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_2_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_2_3_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_2_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_11_), .ZN(
        prince_rounds_SR_Inv_Result_s1[59]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_2_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[10]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_2_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_3_0_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_3_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_12_), .ZN(
        prince_rounds_SR_Inv_Result_s1[12]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_3_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[13]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_3_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_3_1_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_3_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_13_), .ZN(
        prince_rounds_SR_Inv_Result_s1[13]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_3_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s1[13]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_3_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_3_2_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_3_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_14_), .ZN(
        prince_rounds_SR_Inv_Result_s1[14]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_3_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[15]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_3_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_3_3_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_3_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_15_), .ZN(
        prince_rounds_SR_Inv_Result_s1[15]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_3_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[14]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_3_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_4_0_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_4_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_16_), .ZN(
        prince_rounds_SR_Inv_Result_s1[32]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_4_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[17]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_4_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_4_1_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_4_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_17_), .ZN(
        prince_rounds_SR_Inv_Result_s1[33]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_4_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s1[17]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_4_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_4_2_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_4_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_18_), .ZN(
        prince_rounds_SR_Inv_Result_s1[34]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_4_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[19]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_4_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_4_3_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_4_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_19_), .ZN(
        prince_rounds_SR_Inv_Result_s1[35]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_4_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[18]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_4_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_5_0_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_5_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_20_), .ZN(
        prince_rounds_SR_Inv_Result_s1[52]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_5_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[21]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_5_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_5_1_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_5_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_21_), .ZN(
        prince_rounds_SR_Inv_Result_s1[53]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_5_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s1[21]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_5_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_5_2_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_5_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_22_), .ZN(
        prince_rounds_SR_Inv_Result_s1[54]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_5_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[23]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_5_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_5_3_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_5_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_23_), .ZN(
        prince_rounds_SR_Inv_Result_s1[55]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_5_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[22]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_5_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_6_0_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_6_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_24_), .ZN(
        prince_rounds_SR_Inv_Result_s1[8]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_6_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[25]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_6_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_6_1_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_6_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_25_), .ZN(
        prince_rounds_SR_Inv_Result_s1[9]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_6_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s1[25]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_6_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_6_2_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_6_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_26_), .ZN(
        prince_rounds_SR_Inv_Result_s1[10]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_6_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[27]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_6_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_6_3_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_6_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_27_), .ZN(
        prince_rounds_SR_Inv_Result_s1[11]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_6_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[26]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_6_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_7_0_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_7_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_28_), .ZN(
        prince_rounds_SR_Inv_Result_s1[28]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_7_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[29]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_7_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_7_1_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_7_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_29_), .ZN(
        prince_rounds_SR_Inv_Result_s1[29]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_7_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s1[29]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_7_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_7_2_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_7_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_30_), .ZN(
        prince_rounds_SR_Inv_Result_s1[30]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_7_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[31]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_7_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_7_3_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_7_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_31_), .ZN(
        prince_rounds_SR_Inv_Result_s1[31]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_7_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[30]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_7_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_8_0_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_8_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_32_), .ZN(
        prince_rounds_SR_Inv_Result_s1[48]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_8_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[33]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_8_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_8_1_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_8_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_33_), .ZN(
        prince_rounds_SR_Inv_Result_s1[49]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_8_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s1[33]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_8_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_8_2_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_8_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_34_), .ZN(
        prince_rounds_SR_Inv_Result_s1[50]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_8_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[35]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_8_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_8_3_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_8_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_35_), .ZN(
        prince_rounds_SR_Inv_Result_s1[51]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_8_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[34]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_8_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_9_0_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_9_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_36_), .ZN(
        prince_rounds_SR_Inv_Result_s1[4]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_9_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[37]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_9_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_9_1_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_9_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_37_), .ZN(
        prince_rounds_SR_Inv_Result_s1[5]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_9_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s1[37]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_9_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_9_2_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_9_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_38_), .ZN(
        prince_rounds_SR_Inv_Result_s1[6]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_9_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[39]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_9_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_9_3_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_9_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_39_), .ZN(
        prince_rounds_SR_Inv_Result_s1[7]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_9_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[38]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_9_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_10_0_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_10_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_40_), .ZN(
        prince_rounds_SR_Inv_Result_s1[24]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_10_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[41]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_10_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_10_1_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_10_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_41_), .ZN(
        prince_rounds_SR_Inv_Result_s1[25]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_10_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s1[41]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_10_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_10_2_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_10_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_42_), .ZN(
        prince_rounds_SR_Inv_Result_s1[26]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_10_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[43]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_10_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_10_3_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_10_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_43_), .ZN(
        prince_rounds_SR_Inv_Result_s1[27]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_10_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[42]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_10_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_11_0_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_11_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_44_), .ZN(
        prince_rounds_SR_Inv_Result_s1[44]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_11_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[45]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_11_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_11_1_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_11_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_45_), .ZN(
        prince_rounds_SR_Inv_Result_s1[45]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_11_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s1[45]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_11_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_11_2_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_11_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_46_), .ZN(
        prince_rounds_SR_Inv_Result_s1[46]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_11_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[47]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_11_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_11_3_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_11_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_47_), .ZN(
        prince_rounds_SR_Inv_Result_s1[47]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_11_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[46]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_11_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_12_0_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_12_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_48_), .ZN(
        prince_rounds_SR_Inv_Result_s1[0]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_12_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[49]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_12_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_12_1_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_12_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_49_), .ZN(
        prince_rounds_SR_Inv_Result_s1[1]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_12_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s1[49]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_12_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_12_2_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_12_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_50_), .ZN(
        prince_rounds_SR_Inv_Result_s1[2]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_12_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[51]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_12_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_12_3_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_12_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_51_), .ZN(
        prince_rounds_SR_Inv_Result_s1[3]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_12_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[50]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_12_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_13_0_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_13_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_52_), .ZN(
        prince_rounds_SR_Inv_Result_s1[20]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_13_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[53]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_13_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_13_1_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_13_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_53_), .ZN(
        prince_rounds_SR_Inv_Result_s1[21]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_13_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s1[53]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_13_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_13_2_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_13_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_54_), .ZN(
        prince_rounds_SR_Inv_Result_s1[22]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_13_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[55]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_13_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_13_3_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_13_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_55_), .ZN(
        prince_rounds_SR_Inv_Result_s1[23]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_13_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[54]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_13_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_14_0_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_14_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_56_), .ZN(
        prince_rounds_SR_Inv_Result_s1[40]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_14_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[57]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_14_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_14_1_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_14_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_57_), .ZN(
        prince_rounds_SR_Inv_Result_s1[41]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_14_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s1[57]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_14_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_14_2_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_14_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_58_), .ZN(
        prince_rounds_SR_Inv_Result_s1[42]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_14_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[59]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_14_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_14_3_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_14_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_59_), .ZN(
        prince_rounds_SR_Inv_Result_s1[43]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_14_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[58]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_14_3_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_15_0_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_15_0_n3), .B(
        prince_rounds_k1_XOR_round_Constant_60_), .ZN(
        prince_rounds_SR_Inv_Result_s1[60]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_15_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[61]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_15_0_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_15_1_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_15_1_n3), .B(
        prince_rounds_k1_XOR_round_Constant_61_), .ZN(
        prince_rounds_SR_Inv_Result_s1[61]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_15_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s1[61]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_15_1_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_15_2_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_15_2_n3), .B(
        prince_rounds_k1_XOR_round_Constant_62_), .ZN(
        prince_rounds_SR_Inv_Result_s1[62]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_15_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[63]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_15_2_n3) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_15_3_U2 ( .A(
        prince_rounds_AddKey1_forInv_XORInst_15_3_n3), .B(
        prince_rounds_k1_XOR_round_Constant_63_), .ZN(
        prince_rounds_SR_Inv_Result_s1[63]) );
  XNOR2_X1 prince_rounds_AddKey1_forInv_XORInst_15_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s1[62]), .ZN(
        prince_rounds_AddKey1_forInv_XORInst_15_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_0_0_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_0_0_n3), .B(Key2[0]), .ZN(
        prince_rounds_SR_Inv_Result_s2[16]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_0_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[1]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_0_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_0_1_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_0_1_n3), .B(Key2[1]), .ZN(
        prince_rounds_SR_Inv_Result_s2[17]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_0_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s2[1]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_0_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_0_2_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_0_2_n3), .B(Key2[2]), .ZN(
        prince_rounds_SR_Inv_Result_s2[18]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_0_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[3]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_0_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_0_3_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_0_3_n3), .B(Key2[3]), .ZN(
        prince_rounds_SR_Inv_Result_s2[19]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_0_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[2]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_0_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_1_0_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_1_0_n3), .B(Key2[4]), .ZN(
        prince_rounds_SR_Inv_Result_s2[36]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_1_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[5]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_1_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_1_1_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_1_1_n3), .B(Key2[5]), .ZN(
        prince_rounds_SR_Inv_Result_s2[37]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_1_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s2[5]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_1_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_1_2_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_1_2_n3), .B(Key2[6]), .ZN(
        prince_rounds_SR_Inv_Result_s2[38]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_1_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[7]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_1_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_1_3_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_1_3_n3), .B(Key2[7]), .ZN(
        prince_rounds_SR_Inv_Result_s2[39]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_1_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[6]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_1_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_2_0_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_2_0_n3), .B(Key2[8]), .ZN(
        prince_rounds_SR_Inv_Result_s2[56]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_2_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[9]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_2_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_2_1_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_2_1_n3), .B(Key2[9]), .ZN(
        prince_rounds_SR_Inv_Result_s2[57]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_2_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s2[9]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_2_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_2_2_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_2_2_n3), .B(Key2[10]), .ZN(
        prince_rounds_SR_Inv_Result_s2[58]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_2_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[11]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_2_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_2_3_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_2_3_n3), .B(Key2[11]), .ZN(
        prince_rounds_SR_Inv_Result_s2[59]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_2_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[10]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_2_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_3_0_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_3_0_n3), .B(Key2[12]), .ZN(
        prince_rounds_SR_Inv_Result_s2[12]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_3_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[13]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_3_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_3_1_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_3_1_n3), .B(Key2[13]), .ZN(
        prince_rounds_SR_Inv_Result_s2[13]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_3_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s2[13]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_3_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_3_2_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_3_2_n3), .B(Key2[14]), .ZN(
        prince_rounds_SR_Inv_Result_s2[14]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_3_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[15]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_3_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_3_3_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_3_3_n3), .B(Key2[15]), .ZN(
        prince_rounds_SR_Inv_Result_s2[15]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_3_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[14]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_3_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_4_0_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_4_0_n3), .B(Key2[16]), .ZN(
        prince_rounds_SR_Inv_Result_s2[32]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_4_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[17]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_4_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_4_1_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_4_1_n3), .B(Key2[17]), .ZN(
        prince_rounds_SR_Inv_Result_s2[33]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_4_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s2[17]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_4_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_4_2_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_4_2_n3), .B(Key2[18]), .ZN(
        prince_rounds_SR_Inv_Result_s2[34]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_4_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[19]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_4_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_4_3_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_4_3_n3), .B(Key2[19]), .ZN(
        prince_rounds_SR_Inv_Result_s2[35]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_4_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[18]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_4_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_5_0_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_5_0_n3), .B(Key2[20]), .ZN(
        prince_rounds_SR_Inv_Result_s2[52]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_5_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[21]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_5_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_5_1_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_5_1_n3), .B(Key2[21]), .ZN(
        prince_rounds_SR_Inv_Result_s2[53]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_5_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s2[21]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_5_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_5_2_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_5_2_n3), .B(Key2[22]), .ZN(
        prince_rounds_SR_Inv_Result_s2[54]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_5_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[23]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_5_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_5_3_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_5_3_n3), .B(Key2[23]), .ZN(
        prince_rounds_SR_Inv_Result_s2[55]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_5_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[22]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_5_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_6_0_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_6_0_n3), .B(Key2[24]), .ZN(
        prince_rounds_SR_Inv_Result_s2[8]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_6_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[25]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_6_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_6_1_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_6_1_n3), .B(Key2[25]), .ZN(
        prince_rounds_SR_Inv_Result_s2[9]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_6_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s2[25]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_6_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_6_2_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_6_2_n3), .B(Key2[26]), .ZN(
        prince_rounds_SR_Inv_Result_s2[10]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_6_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[27]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_6_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_6_3_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_6_3_n3), .B(Key2[27]), .ZN(
        prince_rounds_SR_Inv_Result_s2[11]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_6_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[26]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_6_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_7_0_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_7_0_n3), .B(Key2[28]), .ZN(
        prince_rounds_SR_Inv_Result_s2[28]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_7_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[29]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_7_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_7_1_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_7_1_n3), .B(Key2[29]), .ZN(
        prince_rounds_SR_Inv_Result_s2[29]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_7_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s2[29]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_7_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_7_2_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_7_2_n3), .B(Key2[30]), .ZN(
        prince_rounds_SR_Inv_Result_s2[30]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_7_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[31]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_7_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_7_3_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_7_3_n3), .B(Key2[31]), .ZN(
        prince_rounds_SR_Inv_Result_s2[31]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_7_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[30]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_7_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_8_0_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_8_0_n3), .B(Key2[32]), .ZN(
        prince_rounds_SR_Inv_Result_s2[48]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_8_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[33]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_8_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_8_1_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_8_1_n3), .B(Key2[33]), .ZN(
        prince_rounds_SR_Inv_Result_s2[49]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_8_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s2[33]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_8_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_8_2_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_8_2_n3), .B(Key2[34]), .ZN(
        prince_rounds_SR_Inv_Result_s2[50]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_8_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[35]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_8_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_8_3_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_8_3_n3), .B(Key2[35]), .ZN(
        prince_rounds_SR_Inv_Result_s2[51]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_8_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[34]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_8_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_9_0_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_9_0_n3), .B(Key2[36]), .ZN(
        prince_rounds_SR_Inv_Result_s2[4]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_9_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[37]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_9_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_9_1_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_9_1_n3), .B(Key2[37]), .ZN(
        prince_rounds_SR_Inv_Result_s2[5]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_9_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s2[37]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_9_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_9_2_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_9_2_n3), .B(Key2[38]), .ZN(
        prince_rounds_SR_Inv_Result_s2[6]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_9_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[39]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_9_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_9_3_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_9_3_n3), .B(Key2[39]), .ZN(
        prince_rounds_SR_Inv_Result_s2[7]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_9_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[38]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_9_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_10_0_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_10_0_n3), .B(Key2[40]), .ZN(
        prince_rounds_SR_Inv_Result_s2[24]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_10_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[41]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_10_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_10_1_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_10_1_n3), .B(Key2[41]), .ZN(
        prince_rounds_SR_Inv_Result_s2[25]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_10_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s2[41]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_10_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_10_2_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_10_2_n3), .B(Key2[42]), .ZN(
        prince_rounds_SR_Inv_Result_s2[26]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_10_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[43]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_10_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_10_3_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_10_3_n3), .B(Key2[43]), .ZN(
        prince_rounds_SR_Inv_Result_s2[27]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_10_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[42]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_10_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_11_0_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_11_0_n3), .B(Key2[44]), .ZN(
        prince_rounds_SR_Inv_Result_s2[44]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_11_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[45]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_11_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_11_1_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_11_1_n3), .B(Key2[45]), .ZN(
        prince_rounds_SR_Inv_Result_s2[45]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_11_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s2[45]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_11_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_11_2_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_11_2_n3), .B(Key2[46]), .ZN(
        prince_rounds_SR_Inv_Result_s2[46]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_11_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[47]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_11_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_11_3_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_11_3_n3), .B(Key2[47]), .ZN(
        prince_rounds_SR_Inv_Result_s2[47]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_11_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[46]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_11_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_12_0_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_12_0_n3), .B(Key2[48]), .ZN(
        prince_rounds_SR_Inv_Result_s2[0]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_12_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[49]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_12_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_12_1_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_12_1_n3), .B(Key2[49]), .ZN(
        prince_rounds_SR_Inv_Result_s2[1]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_12_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s2[49]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_12_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_12_2_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_12_2_n3), .B(Key2[50]), .ZN(
        prince_rounds_SR_Inv_Result_s2[2]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_12_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[51]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_12_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_12_3_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_12_3_n3), .B(Key2[51]), .ZN(
        prince_rounds_SR_Inv_Result_s2[3]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_12_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[50]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_12_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_13_0_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_13_0_n3), .B(Key2[52]), .ZN(
        prince_rounds_SR_Inv_Result_s2[20]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_13_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[53]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_13_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_13_1_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_13_1_n3), .B(Key2[53]), .ZN(
        prince_rounds_SR_Inv_Result_s2[21]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_13_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s2[53]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_13_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_13_2_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_13_2_n3), .B(Key2[54]), .ZN(
        prince_rounds_SR_Inv_Result_s2[22]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_13_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[55]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_13_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_13_3_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_13_3_n3), .B(Key2[55]), .ZN(
        prince_rounds_SR_Inv_Result_s2[23]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_13_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[54]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_13_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_14_0_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_14_0_n3), .B(Key2[56]), .ZN(
        prince_rounds_SR_Inv_Result_s2[40]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_14_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[57]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_14_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_14_1_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_14_1_n3), .B(Key2[57]), .ZN(
        prince_rounds_SR_Inv_Result_s2[41]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_14_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s2[57]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_14_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_14_2_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_14_2_n3), .B(Key2[58]), .ZN(
        prince_rounds_SR_Inv_Result_s2[42]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_14_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[59]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_14_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_14_3_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_14_3_n3), .B(Key2[59]), .ZN(
        prince_rounds_SR_Inv_Result_s2[43]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_14_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[58]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_14_3_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_15_0_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_15_0_n3), .B(Key2[60]), .ZN(
        prince_rounds_SR_Inv_Result_s2[60]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_15_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[61]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_15_0_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_15_1_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_15_1_n3), .B(Key2[61]), .ZN(
        prince_rounds_SR_Inv_Result_s2[61]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_15_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s2[61]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_15_1_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_15_2_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_15_2_n3), .B(Key2[62]), .ZN(
        prince_rounds_SR_Inv_Result_s2[62]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_15_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[63]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_15_2_n3) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_15_3_U2 ( .A(
        prince_rounds_AddKey2_forInv_XORInst_15_3_n3), .B(Key2[63]), .ZN(
        prince_rounds_SR_Inv_Result_s2[63]) );
  XNOR2_X1 prince_rounds_AddKey2_forInv_XORInst_15_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s2[62]), .ZN(
        prince_rounds_AddKey2_forInv_XORInst_15_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_0_0_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_0_0_n3), .B(Key3[0]), .ZN(
        prince_rounds_SR_Inv_Result_s3[16]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_0_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[0]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_0_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_0_1_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_0_1_n3), .B(Key3[1]), .ZN(
        prince_rounds_SR_Inv_Result_s3[17]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_0_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[1]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_0_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_0_2_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_0_2_n3), .B(Key3[2]), .ZN(
        prince_rounds_SR_Inv_Result_s3[18]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_0_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[2]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_0_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_0_3_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_0_3_n3), .B(Key3[3]), .ZN(
        prince_rounds_SR_Inv_Result_s3[19]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_0_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s3[2]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_0_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_1_0_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_1_0_n3), .B(Key3[4]), .ZN(
        prince_rounds_SR_Inv_Result_s3[36]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_1_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[4]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_1_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_1_1_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_1_1_n3), .B(Key3[5]), .ZN(
        prince_rounds_SR_Inv_Result_s3[37]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_1_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[5]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_1_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_1_2_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_1_2_n3), .B(Key3[6]), .ZN(
        prince_rounds_SR_Inv_Result_s3[38]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_1_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[6]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_1_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_1_3_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_1_3_n3), .B(Key3[7]), .ZN(
        prince_rounds_SR_Inv_Result_s3[39]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_1_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s3[6]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_1_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_2_0_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_2_0_n3), .B(Key3[8]), .ZN(
        prince_rounds_SR_Inv_Result_s3[56]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_2_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[8]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_2_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_2_1_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_2_1_n3), .B(Key3[9]), .ZN(
        prince_rounds_SR_Inv_Result_s3[57]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_2_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[9]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_2_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_2_2_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_2_2_n3), .B(Key3[10]), .ZN(
        prince_rounds_SR_Inv_Result_s3[58]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_2_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[10]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_2_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_2_3_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_2_3_n3), .B(Key3[11]), .ZN(
        prince_rounds_SR_Inv_Result_s3[59]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_2_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s3[10]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_2_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_3_0_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_3_0_n3), .B(Key3[12]), .ZN(
        prince_rounds_SR_Inv_Result_s3[12]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_3_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[12]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_3_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_3_1_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_3_1_n3), .B(Key3[13]), .ZN(
        prince_rounds_SR_Inv_Result_s3[13]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_3_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[13]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_3_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_3_2_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_3_2_n3), .B(Key3[14]), .ZN(
        prince_rounds_SR_Inv_Result_s3[14]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_3_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[14]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_3_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_3_3_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_3_3_n3), .B(Key3[15]), .ZN(
        prince_rounds_SR_Inv_Result_s3[15]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_3_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s3[14]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_3_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_4_0_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_4_0_n3), .B(Key3[16]), .ZN(
        prince_rounds_SR_Inv_Result_s3[32]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_4_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[16]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_4_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_4_1_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_4_1_n3), .B(Key3[17]), .ZN(
        prince_rounds_SR_Inv_Result_s3[33]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_4_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[17]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_4_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_4_2_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_4_2_n3), .B(Key3[18]), .ZN(
        prince_rounds_SR_Inv_Result_s3[34]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_4_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[18]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_4_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_4_3_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_4_3_n3), .B(Key3[19]), .ZN(
        prince_rounds_SR_Inv_Result_s3[35]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_4_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s3[18]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_4_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_5_0_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_5_0_n3), .B(Key3[20]), .ZN(
        prince_rounds_SR_Inv_Result_s3[52]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_5_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[20]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_5_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_5_1_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_5_1_n3), .B(Key3[21]), .ZN(
        prince_rounds_SR_Inv_Result_s3[53]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_5_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[21]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_5_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_5_2_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_5_2_n3), .B(Key3[22]), .ZN(
        prince_rounds_SR_Inv_Result_s3[54]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_5_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[22]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_5_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_5_3_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_5_3_n3), .B(Key3[23]), .ZN(
        prince_rounds_SR_Inv_Result_s3[55]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_5_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s3[22]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_5_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_6_0_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_6_0_n3), .B(Key3[24]), .ZN(
        prince_rounds_SR_Inv_Result_s3[8]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_6_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[24]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_6_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_6_1_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_6_1_n3), .B(Key3[25]), .ZN(
        prince_rounds_SR_Inv_Result_s3[9]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_6_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[25]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_6_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_6_2_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_6_2_n3), .B(Key3[26]), .ZN(
        prince_rounds_SR_Inv_Result_s3[10]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_6_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[26]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_6_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_6_3_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_6_3_n3), .B(Key3[27]), .ZN(
        prince_rounds_SR_Inv_Result_s3[11]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_6_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s3[26]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_6_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_7_0_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_7_0_n3), .B(Key3[28]), .ZN(
        prince_rounds_SR_Inv_Result_s3[28]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_7_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[28]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_7_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_7_1_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_7_1_n3), .B(Key3[29]), .ZN(
        prince_rounds_SR_Inv_Result_s3[29]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_7_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[29]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_7_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_7_2_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_7_2_n3), .B(Key3[30]), .ZN(
        prince_rounds_SR_Inv_Result_s3[30]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_7_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[30]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_7_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_7_3_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_7_3_n3), .B(Key3[31]), .ZN(
        prince_rounds_SR_Inv_Result_s3[31]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_7_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s3[30]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_7_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_8_0_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_8_0_n3), .B(Key3[32]), .ZN(
        prince_rounds_SR_Inv_Result_s3[48]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_8_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[32]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_8_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_8_1_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_8_1_n3), .B(Key3[33]), .ZN(
        prince_rounds_SR_Inv_Result_s3[49]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_8_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[33]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_8_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_8_2_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_8_2_n3), .B(Key3[34]), .ZN(
        prince_rounds_SR_Inv_Result_s3[50]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_8_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[34]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_8_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_8_3_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_8_3_n3), .B(Key3[35]), .ZN(
        prince_rounds_SR_Inv_Result_s3[51]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_8_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s3[34]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_8_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_9_0_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_9_0_n3), .B(Key3[36]), .ZN(
        prince_rounds_SR_Inv_Result_s3[4]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_9_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[36]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_9_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_9_1_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_9_1_n3), .B(Key3[37]), .ZN(
        prince_rounds_SR_Inv_Result_s3[5]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_9_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[37]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_9_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_9_2_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_9_2_n3), .B(Key3[38]), .ZN(
        prince_rounds_SR_Inv_Result_s3[6]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_9_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[38]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_9_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_9_3_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_9_3_n3), .B(Key3[39]), .ZN(
        prince_rounds_SR_Inv_Result_s3[7]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_9_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s3[38]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_9_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_10_0_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_10_0_n3), .B(Key3[40]), .ZN(
        prince_rounds_SR_Inv_Result_s3[24]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_10_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[40]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_10_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_10_1_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_10_1_n3), .B(Key3[41]), .ZN(
        prince_rounds_SR_Inv_Result_s3[25]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_10_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[41]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_10_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_10_2_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_10_2_n3), .B(Key3[42]), .ZN(
        prince_rounds_SR_Inv_Result_s3[26]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_10_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[42]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_10_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_10_3_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_10_3_n3), .B(Key3[43]), .ZN(
        prince_rounds_SR_Inv_Result_s3[27]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_10_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s3[42]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_10_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_11_0_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_11_0_n3), .B(Key3[44]), .ZN(
        prince_rounds_SR_Inv_Result_s3[44]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_11_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[44]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_11_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_11_1_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_11_1_n3), .B(Key3[45]), .ZN(
        prince_rounds_SR_Inv_Result_s3[45]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_11_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[45]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_11_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_11_2_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_11_2_n3), .B(Key3[46]), .ZN(
        prince_rounds_SR_Inv_Result_s3[46]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_11_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[46]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_11_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_11_3_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_11_3_n3), .B(Key3[47]), .ZN(
        prince_rounds_SR_Inv_Result_s3[47]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_11_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s3[46]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_11_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_12_0_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_12_0_n3), .B(Key3[48]), .ZN(
        prince_rounds_SR_Inv_Result_s3[0]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_12_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[48]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_12_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_12_1_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_12_1_n3), .B(Key3[49]), .ZN(
        prince_rounds_SR_Inv_Result_s3[1]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_12_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[49]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_12_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_12_2_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_12_2_n3), .B(Key3[50]), .ZN(
        prince_rounds_SR_Inv_Result_s3[2]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_12_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[50]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_12_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_12_3_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_12_3_n3), .B(Key3[51]), .ZN(
        prince_rounds_SR_Inv_Result_s3[3]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_12_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s3[50]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_12_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_13_0_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_13_0_n3), .B(Key3[52]), .ZN(
        prince_rounds_SR_Inv_Result_s3[20]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_13_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[52]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_13_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_13_1_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_13_1_n3), .B(Key3[53]), .ZN(
        prince_rounds_SR_Inv_Result_s3[21]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_13_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[53]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_13_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_13_2_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_13_2_n3), .B(Key3[54]), .ZN(
        prince_rounds_SR_Inv_Result_s3[22]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_13_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[54]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_13_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_13_3_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_13_3_n3), .B(Key3[55]), .ZN(
        prince_rounds_SR_Inv_Result_s3[23]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_13_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s3[54]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_13_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_14_0_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_14_0_n3), .B(Key3[56]), .ZN(
        prince_rounds_SR_Inv_Result_s3[40]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_14_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[56]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_14_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_14_1_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_14_1_n3), .B(Key3[57]), .ZN(
        prince_rounds_SR_Inv_Result_s3[41]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_14_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[57]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_14_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_14_2_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_14_2_n3), .B(Key3[58]), .ZN(
        prince_rounds_SR_Inv_Result_s3[42]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_14_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[58]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_14_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_14_3_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_14_3_n3), .B(Key3[59]), .ZN(
        prince_rounds_SR_Inv_Result_s3[43]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_14_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s3[58]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_14_3_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_15_0_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_15_0_n3), .B(Key3[60]), .ZN(
        prince_rounds_SR_Inv_Result_s3[60]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_15_0_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[60]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_15_0_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_15_1_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_15_1_n3), .B(Key3[61]), .ZN(
        prince_rounds_SR_Inv_Result_s3[61]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_15_1_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[61]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_15_1_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_15_2_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_15_2_n3), .B(Key3[62]), .ZN(
        prince_rounds_SR_Inv_Result_s3[62]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_15_2_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Inv_Result_s3[62]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_15_2_n3) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_15_3_U2 ( .A(
        prince_rounds_AddKey3_forInv_XORInst_15_3_n3), .B(Key3[63]), .ZN(
        prince_rounds_SR_Inv_Result_s3[63]) );
  XNOR2_X1 prince_rounds_AddKey3_forInv_XORInst_15_3_U1 ( .A(1'b0), .B(
        prince_rounds_sub_Result_s3[62]), .ZN(
        prince_rounds_AddKey3_forInv_XORInst_15_3_n3) );
  BUF_X1 prince_rounds_S_Sinv_mul1_U4 ( .A(roundEnd_Select_Signal), .Z(
        prince_rounds_S_Sinv_mul1_n8) );
  BUF_X1 prince_rounds_S_Sinv_mul1_U3 ( .A(prince_rounds_S_Sinv_mul1_n8), .Z(
        prince_rounds_S_Sinv_mul1_n10) );
  BUF_X1 prince_rounds_S_Sinv_mul1_U2 ( .A(roundEnd_Select_Signal), .Z(
        prince_rounds_S_Sinv_mul1_n7) );
  BUF_X1 prince_rounds_S_Sinv_mul1_U1 ( .A(prince_rounds_S_Sinv_mul1_n7), .Z(
        prince_rounds_S_Sinv_mul1_n9) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_0_U1 ( .A(
        prince_rounds_sub_Result_s1[0]), .B(prince_rounds_SR_Inv_Result_s1[0]), 
        .S(prince_rounds_S_Sinv_mul1_n9), .Z(prince_rounds_mul_input_s1[0]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_1_U1 ( .A(
        prince_rounds_sub_Result_s1[1]), .B(prince_rounds_SR_Inv_Result_s1[1]), 
        .S(prince_rounds_S_Sinv_mul1_n9), .Z(prince_rounds_mul_input_s1[1]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_2_U1 ( .A(
        prince_rounds_sub_Result_s1[2]), .B(prince_rounds_SR_Inv_Result_s1[2]), 
        .S(prince_rounds_S_Sinv_mul1_n9), .Z(prince_rounds_mul_input_s1[2]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_3_U1 ( .A(
        prince_rounds_sub_Result_s1[3]), .B(prince_rounds_SR_Inv_Result_s1[3]), 
        .S(prince_rounds_S_Sinv_mul1_n9), .Z(prince_rounds_mul_input_s1[3]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_4_U1 ( .A(
        prince_rounds_sub_Result_s1[4]), .B(prince_rounds_SR_Inv_Result_s1[4]), 
        .S(prince_rounds_S_Sinv_mul1_n9), .Z(prince_rounds_mul_input_s1[4]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_5_U1 ( .A(
        prince_rounds_sub_Result_s1[5]), .B(prince_rounds_SR_Inv_Result_s1[5]), 
        .S(prince_rounds_S_Sinv_mul1_n9), .Z(prince_rounds_mul_input_s1[5]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_6_U1 ( .A(
        prince_rounds_sub_Result_s1[6]), .B(prince_rounds_SR_Inv_Result_s1[6]), 
        .S(prince_rounds_S_Sinv_mul1_n9), .Z(prince_rounds_mul_input_s1[6]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_7_U1 ( .A(
        prince_rounds_sub_Result_s1[7]), .B(prince_rounds_SR_Inv_Result_s1[7]), 
        .S(prince_rounds_S_Sinv_mul1_n9), .Z(prince_rounds_mul_input_s1[7]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_8_U1 ( .A(
        prince_rounds_sub_Result_s1[8]), .B(prince_rounds_SR_Inv_Result_s1[8]), 
        .S(prince_rounds_S_Sinv_mul1_n9), .Z(prince_rounds_mul_input_s1[8]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_9_U1 ( .A(
        prince_rounds_sub_Result_s1[9]), .B(prince_rounds_SR_Inv_Result_s1[9]), 
        .S(prince_rounds_S_Sinv_mul1_n9), .Z(prince_rounds_mul_input_s1[9]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_10_U1 ( .A(
        prince_rounds_sub_Result_s1[10]), .B(
        prince_rounds_SR_Inv_Result_s1[10]), .S(prince_rounds_S_Sinv_mul1_n9), 
        .Z(prince_rounds_mul_input_s1[10]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_11_U1 ( .A(
        prince_rounds_sub_Result_s1[11]), .B(
        prince_rounds_SR_Inv_Result_s1[11]), .S(prince_rounds_S_Sinv_mul1_n9), 
        .Z(prince_rounds_mul_input_s1[11]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_12_U1 ( .A(
        prince_rounds_sub_Result_s1[12]), .B(
        prince_rounds_SR_Inv_Result_s1[12]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[12]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_13_U1 ( .A(
        prince_rounds_sub_Result_s1[13]), .B(
        prince_rounds_SR_Inv_Result_s1[13]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[13]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_14_U1 ( .A(
        prince_rounds_sub_Result_s1[14]), .B(
        prince_rounds_SR_Inv_Result_s1[14]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[14]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_15_U1 ( .A(
        prince_rounds_sub_Result_s1[15]), .B(
        prince_rounds_SR_Inv_Result_s1[15]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[15]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_16_U1 ( .A(
        prince_rounds_sub_Result_s1[16]), .B(
        prince_rounds_SR_Inv_Result_s1[16]), .S(prince_rounds_S_Sinv_mul1_n9), 
        .Z(prince_rounds_mul_input_s1[16]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_17_U1 ( .A(
        prince_rounds_sub_Result_s1[17]), .B(
        prince_rounds_SR_Inv_Result_s1[17]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[17]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_18_U1 ( .A(
        prince_rounds_sub_Result_s1[18]), .B(
        prince_rounds_SR_Inv_Result_s1[18]), .S(prince_rounds_S_Sinv_mul1_n9), 
        .Z(prince_rounds_mul_input_s1[18]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_19_U1 ( .A(
        prince_rounds_sub_Result_s1[19]), .B(
        prince_rounds_SR_Inv_Result_s1[19]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[19]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_20_U1 ( .A(
        prince_rounds_sub_Result_s1[20]), .B(
        prince_rounds_SR_Inv_Result_s1[20]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[20]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_21_U1 ( .A(
        prince_rounds_sub_Result_s1[21]), .B(
        prince_rounds_SR_Inv_Result_s1[21]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[21]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_22_U1 ( .A(
        prince_rounds_sub_Result_s1[22]), .B(
        prince_rounds_SR_Inv_Result_s1[22]), .S(prince_rounds_S_Sinv_mul1_n9), 
        .Z(prince_rounds_mul_input_s1[22]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_23_U1 ( .A(
        prince_rounds_sub_Result_s1[23]), .B(
        prince_rounds_SR_Inv_Result_s1[23]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[23]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_24_U1 ( .A(
        prince_rounds_sub_Result_s1[24]), .B(
        prince_rounds_SR_Inv_Result_s1[24]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[24]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_25_U1 ( .A(
        prince_rounds_sub_Result_s1[25]), .B(
        prince_rounds_SR_Inv_Result_s1[25]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[25]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_26_U1 ( .A(
        prince_rounds_sub_Result_s1[26]), .B(
        prince_rounds_SR_Inv_Result_s1[26]), .S(prince_rounds_S_Sinv_mul1_n9), 
        .Z(prince_rounds_mul_input_s1[26]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_27_U1 ( .A(
        prince_rounds_sub_Result_s1[27]), .B(
        prince_rounds_SR_Inv_Result_s1[27]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[27]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_28_U1 ( .A(
        prince_rounds_sub_Result_s1[28]), .B(
        prince_rounds_SR_Inv_Result_s1[28]), .S(prince_rounds_S_Sinv_mul1_n9), 
        .Z(prince_rounds_mul_input_s1[28]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_29_U1 ( .A(
        prince_rounds_sub_Result_s1[29]), .B(
        prince_rounds_SR_Inv_Result_s1[29]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[29]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_30_U1 ( .A(
        prince_rounds_sub_Result_s1[30]), .B(
        prince_rounds_SR_Inv_Result_s1[30]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[30]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_31_U1 ( .A(
        prince_rounds_sub_Result_s1[31]), .B(
        prince_rounds_SR_Inv_Result_s1[31]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[31]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_32_U1 ( .A(
        prince_rounds_sub_Result_s1[32]), .B(
        prince_rounds_SR_Inv_Result_s1[32]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[32]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_33_U1 ( .A(
        prince_rounds_sub_Result_s1[33]), .B(
        prince_rounds_SR_Inv_Result_s1[33]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[33]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_34_U1 ( .A(
        prince_rounds_sub_Result_s1[34]), .B(
        prince_rounds_SR_Inv_Result_s1[34]), .S(prince_rounds_S_Sinv_mul1_n9), 
        .Z(prince_rounds_mul_input_s1[34]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_35_U1 ( .A(
        prince_rounds_sub_Result_s1[35]), .B(
        prince_rounds_SR_Inv_Result_s1[35]), .S(prince_rounds_S_Sinv_mul1_n7), 
        .Z(prince_rounds_mul_input_s1[35]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_36_U1 ( .A(
        prince_rounds_sub_Result_s1[36]), .B(
        prince_rounds_SR_Inv_Result_s1[36]), .S(prince_rounds_S_Sinv_mul1_n10), 
        .Z(prince_rounds_mul_input_s1[36]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_37_U1 ( .A(
        prince_rounds_sub_Result_s1[37]), .B(
        prince_rounds_SR_Inv_Result_s1[37]), .S(prince_rounds_S_Sinv_mul1_n10), 
        .Z(prince_rounds_mul_input_s1[37]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_38_U1 ( .A(
        prince_rounds_sub_Result_s1[38]), .B(
        prince_rounds_SR_Inv_Result_s1[38]), .S(prince_rounds_S_Sinv_mul1_n10), 
        .Z(prince_rounds_mul_input_s1[38]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_39_U1 ( .A(
        prince_rounds_sub_Result_s1[39]), .B(
        prince_rounds_SR_Inv_Result_s1[39]), .S(prince_rounds_S_Sinv_mul1_n10), 
        .Z(prince_rounds_mul_input_s1[39]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_40_U1 ( .A(
        prince_rounds_sub_Result_s1[40]), .B(
        prince_rounds_SR_Inv_Result_s1[40]), .S(prince_rounds_S_Sinv_mul1_n10), 
        .Z(prince_rounds_mul_input_s1[40]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_41_U1 ( .A(
        prince_rounds_sub_Result_s1[41]), .B(
        prince_rounds_SR_Inv_Result_s1[41]), .S(prince_rounds_S_Sinv_mul1_n10), 
        .Z(prince_rounds_mul_input_s1[41]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_42_U1 ( .A(
        prince_rounds_sub_Result_s1[42]), .B(
        prince_rounds_SR_Inv_Result_s1[42]), .S(prince_rounds_S_Sinv_mul1_n10), 
        .Z(prince_rounds_mul_input_s1[42]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_43_U1 ( .A(
        prince_rounds_sub_Result_s1[43]), .B(
        prince_rounds_SR_Inv_Result_s1[43]), .S(prince_rounds_S_Sinv_mul1_n10), 
        .Z(prince_rounds_mul_input_s1[43]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_44_U1 ( .A(
        prince_rounds_sub_Result_s1[44]), .B(
        prince_rounds_SR_Inv_Result_s1[44]), .S(prince_rounds_S_Sinv_mul1_n10), 
        .Z(prince_rounds_mul_input_s1[44]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_45_U1 ( .A(
        prince_rounds_sub_Result_s1[45]), .B(
        prince_rounds_SR_Inv_Result_s1[45]), .S(prince_rounds_S_Sinv_mul1_n10), 
        .Z(prince_rounds_mul_input_s1[45]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_46_U1 ( .A(
        prince_rounds_sub_Result_s1[46]), .B(
        prince_rounds_SR_Inv_Result_s1[46]), .S(prince_rounds_S_Sinv_mul1_n10), 
        .Z(prince_rounds_mul_input_s1[46]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_47_U1 ( .A(
        prince_rounds_sub_Result_s1[47]), .B(
        prince_rounds_SR_Inv_Result_s1[47]), .S(prince_rounds_S_Sinv_mul1_n10), 
        .Z(prince_rounds_mul_input_s1[47]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_48_U1 ( .A(
        prince_rounds_sub_Result_s1[48]), .B(
        prince_rounds_SR_Inv_Result_s1[48]), .S(prince_rounds_S_Sinv_mul1_n10), 
        .Z(prince_rounds_mul_input_s1[48]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_49_U1 ( .A(
        prince_rounds_sub_Result_s1[49]), .B(
        prince_rounds_SR_Inv_Result_s1[49]), .S(prince_rounds_S_Sinv_mul1_n8), 
        .Z(prince_rounds_mul_input_s1[49]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_50_U1 ( .A(
        prince_rounds_sub_Result_s1[50]), .B(
        prince_rounds_SR_Inv_Result_s1[50]), .S(prince_rounds_S_Sinv_mul1_n8), 
        .Z(prince_rounds_mul_input_s1[50]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_51_U1 ( .A(
        prince_rounds_sub_Result_s1[51]), .B(
        prince_rounds_SR_Inv_Result_s1[51]), .S(prince_rounds_S_Sinv_mul1_n8), 
        .Z(prince_rounds_mul_input_s1[51]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_52_U1 ( .A(
        prince_rounds_sub_Result_s1[52]), .B(
        prince_rounds_SR_Inv_Result_s1[52]), .S(prince_rounds_S_Sinv_mul1_n8), 
        .Z(prince_rounds_mul_input_s1[52]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_53_U1 ( .A(
        prince_rounds_sub_Result_s1[53]), .B(
        prince_rounds_SR_Inv_Result_s1[53]), .S(prince_rounds_S_Sinv_mul1_n8), 
        .Z(prince_rounds_mul_input_s1[53]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_54_U1 ( .A(
        prince_rounds_sub_Result_s1[54]), .B(
        prince_rounds_SR_Inv_Result_s1[54]), .S(prince_rounds_S_Sinv_mul1_n8), 
        .Z(prince_rounds_mul_input_s1[54]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_55_U1 ( .A(
        prince_rounds_sub_Result_s1[55]), .B(
        prince_rounds_SR_Inv_Result_s1[55]), .S(prince_rounds_S_Sinv_mul1_n8), 
        .Z(prince_rounds_mul_input_s1[55]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_56_U1 ( .A(
        prince_rounds_sub_Result_s1[56]), .B(
        prince_rounds_SR_Inv_Result_s1[56]), .S(prince_rounds_S_Sinv_mul1_n8), 
        .Z(prince_rounds_mul_input_s1[56]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_57_U1 ( .A(
        prince_rounds_sub_Result_s1[57]), .B(
        prince_rounds_SR_Inv_Result_s1[57]), .S(prince_rounds_S_Sinv_mul1_n8), 
        .Z(prince_rounds_mul_input_s1[57]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_58_U1 ( .A(
        prince_rounds_sub_Result_s1[58]), .B(
        prince_rounds_SR_Inv_Result_s1[58]), .S(prince_rounds_S_Sinv_mul1_n8), 
        .Z(prince_rounds_mul_input_s1[58]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_59_U1 ( .A(
        prince_rounds_sub_Result_s1[59]), .B(
        prince_rounds_SR_Inv_Result_s1[59]), .S(prince_rounds_S_Sinv_mul1_n8), 
        .Z(prince_rounds_mul_input_s1[59]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_60_U1 ( .A(
        prince_rounds_sub_Result_s1[60]), .B(
        prince_rounds_SR_Inv_Result_s1[60]), .S(prince_rounds_S_Sinv_mul1_n10), 
        .Z(prince_rounds_mul_input_s1[60]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_61_U1 ( .A(
        prince_rounds_sub_Result_s1[61]), .B(
        prince_rounds_SR_Inv_Result_s1[61]), .S(prince_rounds_S_Sinv_mul1_n8), 
        .Z(prince_rounds_mul_input_s1[61]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_62_U1 ( .A(
        prince_rounds_sub_Result_s1[62]), .B(
        prince_rounds_SR_Inv_Result_s1[62]), .S(prince_rounds_S_Sinv_mul1_n8), 
        .Z(prince_rounds_mul_input_s1[62]) );
  MUX2_X1 prince_rounds_S_Sinv_mul1_MUXInst_63_U1 ( .A(
        prince_rounds_sub_Result_s1[63]), .B(
        prince_rounds_SR_Inv_Result_s1[63]), .S(prince_rounds_S_Sinv_mul1_n8), 
        .Z(prince_rounds_mul_input_s1[63]) );
  BUF_X1 prince_rounds_S_Sinv_mul2_U4 ( .A(roundEnd_Select_Signal), .Z(
        prince_rounds_S_Sinv_mul2_n7) );
  BUF_X1 prince_rounds_S_Sinv_mul2_U3 ( .A(prince_rounds_S_Sinv_mul2_n7), .Z(
        prince_rounds_S_Sinv_mul2_n9) );
  BUF_X1 prince_rounds_S_Sinv_mul2_U2 ( .A(roundEnd_Select_Signal), .Z(
        prince_rounds_S_Sinv_mul2_n8) );
  BUF_X1 prince_rounds_S_Sinv_mul2_U1 ( .A(prince_rounds_S_Sinv_mul2_n8), .Z(
        prince_rounds_S_Sinv_mul2_n10) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_0_U1 ( .A(
        prince_rounds_sub_Result_s2[0]), .B(prince_rounds_SR_Inv_Result_s2[0]), 
        .S(prince_rounds_S_Sinv_mul2_n9), .Z(prince_rounds_mul_input_s2[0]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_1_U1 ( .A(
        prince_rounds_sub_Result_s2[1]), .B(prince_rounds_SR_Inv_Result_s2[1]), 
        .S(prince_rounds_S_Sinv_mul2_n9), .Z(prince_rounds_mul_input_s2[1]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_2_U1 ( .A(
        prince_rounds_sub_Result_s2[2]), .B(prince_rounds_SR_Inv_Result_s2[2]), 
        .S(prince_rounds_S_Sinv_mul2_n9), .Z(prince_rounds_mul_input_s2[2]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_3_U1 ( .A(
        prince_rounds_sub_Result_s2[3]), .B(prince_rounds_SR_Inv_Result_s2[3]), 
        .S(prince_rounds_S_Sinv_mul2_n9), .Z(prince_rounds_mul_input_s2[3]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_4_U1 ( .A(
        prince_rounds_sub_Result_s2[4]), .B(prince_rounds_SR_Inv_Result_s2[4]), 
        .S(prince_rounds_S_Sinv_mul2_n9), .Z(prince_rounds_mul_input_s2[4]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_5_U1 ( .A(
        prince_rounds_sub_Result_s2[5]), .B(prince_rounds_SR_Inv_Result_s2[5]), 
        .S(prince_rounds_S_Sinv_mul2_n9), .Z(prince_rounds_mul_input_s2[5]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_6_U1 ( .A(
        prince_rounds_sub_Result_s2[6]), .B(prince_rounds_SR_Inv_Result_s2[6]), 
        .S(prince_rounds_S_Sinv_mul2_n9), .Z(prince_rounds_mul_input_s2[6]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_7_U1 ( .A(
        prince_rounds_sub_Result_s2[7]), .B(prince_rounds_SR_Inv_Result_s2[7]), 
        .S(prince_rounds_S_Sinv_mul2_n9), .Z(prince_rounds_mul_input_s2[7]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_8_U1 ( .A(
        prince_rounds_sub_Result_s2[8]), .B(prince_rounds_SR_Inv_Result_s2[8]), 
        .S(prince_rounds_S_Sinv_mul2_n9), .Z(prince_rounds_mul_input_s2[8]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_9_U1 ( .A(
        prince_rounds_sub_Result_s2[9]), .B(prince_rounds_SR_Inv_Result_s2[9]), 
        .S(prince_rounds_S_Sinv_mul2_n9), .Z(prince_rounds_mul_input_s2[9]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_10_U1 ( .A(
        prince_rounds_sub_Result_s2[10]), .B(
        prince_rounds_SR_Inv_Result_s2[10]), .S(prince_rounds_S_Sinv_mul2_n9), 
        .Z(prince_rounds_mul_input_s2[10]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_11_U1 ( .A(
        prince_rounds_sub_Result_s2[11]), .B(
        prince_rounds_SR_Inv_Result_s2[11]), .S(prince_rounds_S_Sinv_mul2_n9), 
        .Z(prince_rounds_mul_input_s2[11]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_12_U1 ( .A(
        prince_rounds_sub_Result_s2[12]), .B(
        prince_rounds_SR_Inv_Result_s2[12]), .S(prince_rounds_S_Sinv_mul2_n9), 
        .Z(prince_rounds_mul_input_s2[12]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_13_U1 ( .A(
        prince_rounds_sub_Result_s2[13]), .B(
        prince_rounds_SR_Inv_Result_s2[13]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[13]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_14_U1 ( .A(
        prince_rounds_sub_Result_s2[14]), .B(
        prince_rounds_SR_Inv_Result_s2[14]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[14]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_15_U1 ( .A(
        prince_rounds_sub_Result_s2[15]), .B(
        prince_rounds_SR_Inv_Result_s2[15]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[15]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_16_U1 ( .A(
        prince_rounds_sub_Result_s2[16]), .B(
        prince_rounds_SR_Inv_Result_s2[16]), .S(prince_rounds_S_Sinv_mul2_n9), 
        .Z(prince_rounds_mul_input_s2[16]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_17_U1 ( .A(
        prince_rounds_sub_Result_s2[17]), .B(
        prince_rounds_SR_Inv_Result_s2[17]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[17]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_18_U1 ( .A(
        prince_rounds_sub_Result_s2[18]), .B(
        prince_rounds_SR_Inv_Result_s2[18]), .S(prince_rounds_S_Sinv_mul2_n9), 
        .Z(prince_rounds_mul_input_s2[18]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_19_U1 ( .A(
        prince_rounds_sub_Result_s2[19]), .B(
        prince_rounds_SR_Inv_Result_s2[19]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[19]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_20_U1 ( .A(
        prince_rounds_sub_Result_s2[20]), .B(
        prince_rounds_SR_Inv_Result_s2[20]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[20]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_21_U1 ( .A(
        prince_rounds_sub_Result_s2[21]), .B(
        prince_rounds_SR_Inv_Result_s2[21]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[21]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_22_U1 ( .A(
        prince_rounds_sub_Result_s2[22]), .B(
        prince_rounds_SR_Inv_Result_s2[22]), .S(prince_rounds_S_Sinv_mul2_n9), 
        .Z(prince_rounds_mul_input_s2[22]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_23_U1 ( .A(
        prince_rounds_sub_Result_s2[23]), .B(
        prince_rounds_SR_Inv_Result_s2[23]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[23]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_24_U1 ( .A(
        prince_rounds_sub_Result_s2[24]), .B(
        prince_rounds_SR_Inv_Result_s2[24]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[24]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_25_U1 ( .A(
        prince_rounds_sub_Result_s2[25]), .B(
        prince_rounds_SR_Inv_Result_s2[25]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[25]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_26_U1 ( .A(
        prince_rounds_sub_Result_s2[26]), .B(
        prince_rounds_SR_Inv_Result_s2[26]), .S(prince_rounds_S_Sinv_mul2_n9), 
        .Z(prince_rounds_mul_input_s2[26]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_27_U1 ( .A(
        prince_rounds_sub_Result_s2[27]), .B(
        prince_rounds_SR_Inv_Result_s2[27]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[27]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_28_U1 ( .A(
        prince_rounds_sub_Result_s2[28]), .B(
        prince_rounds_SR_Inv_Result_s2[28]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[28]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_29_U1 ( .A(
        prince_rounds_sub_Result_s2[29]), .B(
        prince_rounds_SR_Inv_Result_s2[29]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[29]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_30_U1 ( .A(
        prince_rounds_sub_Result_s2[30]), .B(
        prince_rounds_SR_Inv_Result_s2[30]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[30]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_31_U1 ( .A(
        prince_rounds_sub_Result_s2[31]), .B(
        prince_rounds_SR_Inv_Result_s2[31]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[31]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_32_U1 ( .A(
        prince_rounds_sub_Result_s2[32]), .B(
        prince_rounds_SR_Inv_Result_s2[32]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[32]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_33_U1 ( .A(
        prince_rounds_sub_Result_s2[33]), .B(
        prince_rounds_SR_Inv_Result_s2[33]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[33]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_34_U1 ( .A(
        prince_rounds_sub_Result_s2[34]), .B(
        prince_rounds_SR_Inv_Result_s2[34]), .S(prince_rounds_S_Sinv_mul2_n9), 
        .Z(prince_rounds_mul_input_s2[34]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_35_U1 ( .A(
        prince_rounds_sub_Result_s2[35]), .B(
        prince_rounds_SR_Inv_Result_s2[35]), .S(prince_rounds_S_Sinv_mul2_n7), 
        .Z(prince_rounds_mul_input_s2[35]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_36_U1 ( .A(
        prince_rounds_sub_Result_s2[36]), .B(
        prince_rounds_SR_Inv_Result_s2[36]), .S(prince_rounds_S_Sinv_mul2_n10), 
        .Z(prince_rounds_mul_input_s2[36]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_37_U1 ( .A(
        prince_rounds_sub_Result_s2[37]), .B(
        prince_rounds_SR_Inv_Result_s2[37]), .S(prince_rounds_S_Sinv_mul2_n10), 
        .Z(prince_rounds_mul_input_s2[37]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_38_U1 ( .A(
        prince_rounds_sub_Result_s2[38]), .B(
        prince_rounds_SR_Inv_Result_s2[38]), .S(prince_rounds_S_Sinv_mul2_n10), 
        .Z(prince_rounds_mul_input_s2[38]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_39_U1 ( .A(
        prince_rounds_sub_Result_s2[39]), .B(
        prince_rounds_SR_Inv_Result_s2[39]), .S(prince_rounds_S_Sinv_mul2_n10), 
        .Z(prince_rounds_mul_input_s2[39]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_40_U1 ( .A(
        prince_rounds_sub_Result_s2[40]), .B(
        prince_rounds_SR_Inv_Result_s2[40]), .S(prince_rounds_S_Sinv_mul2_n10), 
        .Z(prince_rounds_mul_input_s2[40]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_41_U1 ( .A(
        prince_rounds_sub_Result_s2[41]), .B(
        prince_rounds_SR_Inv_Result_s2[41]), .S(prince_rounds_S_Sinv_mul2_n10), 
        .Z(prince_rounds_mul_input_s2[41]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_42_U1 ( .A(
        prince_rounds_sub_Result_s2[42]), .B(
        prince_rounds_SR_Inv_Result_s2[42]), .S(prince_rounds_S_Sinv_mul2_n10), 
        .Z(prince_rounds_mul_input_s2[42]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_43_U1 ( .A(
        prince_rounds_sub_Result_s2[43]), .B(
        prince_rounds_SR_Inv_Result_s2[43]), .S(prince_rounds_S_Sinv_mul2_n10), 
        .Z(prince_rounds_mul_input_s2[43]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_44_U1 ( .A(
        prince_rounds_sub_Result_s2[44]), .B(
        prince_rounds_SR_Inv_Result_s2[44]), .S(prince_rounds_S_Sinv_mul2_n10), 
        .Z(prince_rounds_mul_input_s2[44]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_45_U1 ( .A(
        prince_rounds_sub_Result_s2[45]), .B(
        prince_rounds_SR_Inv_Result_s2[45]), .S(prince_rounds_S_Sinv_mul2_n10), 
        .Z(prince_rounds_mul_input_s2[45]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_46_U1 ( .A(
        prince_rounds_sub_Result_s2[46]), .B(
        prince_rounds_SR_Inv_Result_s2[46]), .S(prince_rounds_S_Sinv_mul2_n10), 
        .Z(prince_rounds_mul_input_s2[46]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_47_U1 ( .A(
        prince_rounds_sub_Result_s2[47]), .B(
        prince_rounds_SR_Inv_Result_s2[47]), .S(prince_rounds_S_Sinv_mul2_n10), 
        .Z(prince_rounds_mul_input_s2[47]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_48_U1 ( .A(
        prince_rounds_sub_Result_s2[48]), .B(
        prince_rounds_SR_Inv_Result_s2[48]), .S(prince_rounds_S_Sinv_mul2_n10), 
        .Z(prince_rounds_mul_input_s2[48]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_49_U1 ( .A(
        prince_rounds_sub_Result_s2[49]), .B(
        prince_rounds_SR_Inv_Result_s2[49]), .S(prince_rounds_S_Sinv_mul2_n8), 
        .Z(prince_rounds_mul_input_s2[49]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_50_U1 ( .A(
        prince_rounds_sub_Result_s2[50]), .B(
        prince_rounds_SR_Inv_Result_s2[50]), .S(prince_rounds_S_Sinv_mul2_n8), 
        .Z(prince_rounds_mul_input_s2[50]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_51_U1 ( .A(
        prince_rounds_sub_Result_s2[51]), .B(
        prince_rounds_SR_Inv_Result_s2[51]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s2[51]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_52_U1 ( .A(
        prince_rounds_sub_Result_s2[52]), .B(
        prince_rounds_SR_Inv_Result_s2[52]), .S(prince_rounds_S_Sinv_mul2_n8), 
        .Z(prince_rounds_mul_input_s2[52]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_53_U1 ( .A(
        prince_rounds_sub_Result_s2[53]), .B(
        prince_rounds_SR_Inv_Result_s2[53]), .S(prince_rounds_S_Sinv_mul2_n8), 
        .Z(prince_rounds_mul_input_s2[53]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_54_U1 ( .A(
        prince_rounds_sub_Result_s2[54]), .B(
        prince_rounds_SR_Inv_Result_s2[54]), .S(prince_rounds_S_Sinv_mul2_n8), 
        .Z(prince_rounds_mul_input_s2[54]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_55_U1 ( .A(
        prince_rounds_sub_Result_s2[55]), .B(
        prince_rounds_SR_Inv_Result_s2[55]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s2[55]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_56_U1 ( .A(
        prince_rounds_sub_Result_s2[56]), .B(
        prince_rounds_SR_Inv_Result_s2[56]), .S(prince_rounds_S_Sinv_mul2_n8), 
        .Z(prince_rounds_mul_input_s2[56]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_57_U1 ( .A(
        prince_rounds_sub_Result_s2[57]), .B(
        prince_rounds_SR_Inv_Result_s2[57]), .S(prince_rounds_S_Sinv_mul2_n8), 
        .Z(prince_rounds_mul_input_s2[57]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_58_U1 ( .A(
        prince_rounds_sub_Result_s2[58]), .B(
        prince_rounds_SR_Inv_Result_s2[58]), .S(prince_rounds_S_Sinv_mul2_n8), 
        .Z(prince_rounds_mul_input_s2[58]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_59_U1 ( .A(
        prince_rounds_sub_Result_s2[59]), .B(
        prince_rounds_SR_Inv_Result_s2[59]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s2[59]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_60_U1 ( .A(
        prince_rounds_sub_Result_s2[60]), .B(
        prince_rounds_SR_Inv_Result_s2[60]), .S(prince_rounds_S_Sinv_mul2_n10), 
        .Z(prince_rounds_mul_input_s2[60]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_61_U1 ( .A(
        prince_rounds_sub_Result_s2[61]), .B(
        prince_rounds_SR_Inv_Result_s2[61]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s2[61]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_62_U1 ( .A(
        prince_rounds_sub_Result_s2[62]), .B(
        prince_rounds_SR_Inv_Result_s2[62]), .S(prince_rounds_S_Sinv_mul2_n8), 
        .Z(prince_rounds_mul_input_s2[62]) );
  MUX2_X1 prince_rounds_S_Sinv_mul2_MUXInst_63_U1 ( .A(
        prince_rounds_sub_Result_s2[63]), .B(
        prince_rounds_SR_Inv_Result_s2[63]), .S(prince_rounds_S_Sinv_mul2_n8), 
        .Z(prince_rounds_mul_input_s2[63]) );
  BUF_X1 prince_rounds_S_Sinv_mul3_U3 ( .A(roundEnd_Select_Signal), .Z(
        prince_rounds_S_Sinv_mul3_n6) );
  BUF_X1 prince_rounds_S_Sinv_mul3_U2 ( .A(prince_rounds_S_Sinv_mul3_n6), .Z(
        prince_rounds_S_Sinv_mul3_n8) );
  BUF_X1 prince_rounds_S_Sinv_mul3_U1 ( .A(roundEnd_Select_Signal), .Z(
        prince_rounds_S_Sinv_mul3_n7) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_0_U1 ( .A(
        prince_rounds_sub_Result_s3[0]), .B(prince_rounds_SR_Inv_Result_s3[0]), 
        .S(prince_rounds_S_Sinv_mul3_n8), .Z(prince_rounds_mul_input_s3[0]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_1_U1 ( .A(
        prince_rounds_sub_Result_s3[1]), .B(prince_rounds_SR_Inv_Result_s3[1]), 
        .S(prince_rounds_S_Sinv_mul3_n8), .Z(prince_rounds_mul_input_s3[1]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_2_U1 ( .A(
        prince_rounds_sub_Result_s3[2]), .B(prince_rounds_SR_Inv_Result_s3[2]), 
        .S(prince_rounds_S_Sinv_mul3_n8), .Z(prince_rounds_mul_input_s3[2]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_3_U1 ( .A(
        prince_rounds_sub_Result_s3[3]), .B(prince_rounds_SR_Inv_Result_s3[3]), 
        .S(prince_rounds_S_Sinv_mul3_n8), .Z(prince_rounds_mul_input_s3[3]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_4_U1 ( .A(
        prince_rounds_sub_Result_s3[4]), .B(prince_rounds_SR_Inv_Result_s3[4]), 
        .S(prince_rounds_S_Sinv_mul3_n8), .Z(prince_rounds_mul_input_s3[4]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_5_U1 ( .A(
        prince_rounds_sub_Result_s3[5]), .B(prince_rounds_SR_Inv_Result_s3[5]), 
        .S(prince_rounds_S_Sinv_mul3_n8), .Z(prince_rounds_mul_input_s3[5]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_6_U1 ( .A(
        prince_rounds_sub_Result_s3[6]), .B(prince_rounds_SR_Inv_Result_s3[6]), 
        .S(prince_rounds_S_Sinv_mul3_n8), .Z(prince_rounds_mul_input_s3[6]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_7_U1 ( .A(
        prince_rounds_sub_Result_s3[7]), .B(prince_rounds_SR_Inv_Result_s3[7]), 
        .S(prince_rounds_S_Sinv_mul3_n8), .Z(prince_rounds_mul_input_s3[7]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_8_U1 ( .A(
        prince_rounds_sub_Result_s3[8]), .B(prince_rounds_SR_Inv_Result_s3[8]), 
        .S(prince_rounds_S_Sinv_mul3_n8), .Z(prince_rounds_mul_input_s3[8]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_9_U1 ( .A(
        prince_rounds_sub_Result_s3[9]), .B(prince_rounds_SR_Inv_Result_s3[9]), 
        .S(prince_rounds_S_Sinv_mul3_n8), .Z(prince_rounds_mul_input_s3[9]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_10_U1 ( .A(
        prince_rounds_sub_Result_s3[10]), .B(
        prince_rounds_SR_Inv_Result_s3[10]), .S(prince_rounds_S_Sinv_mul3_n8), 
        .Z(prince_rounds_mul_input_s3[10]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_11_U1 ( .A(
        prince_rounds_sub_Result_s3[11]), .B(
        prince_rounds_SR_Inv_Result_s3[11]), .S(prince_rounds_S_Sinv_mul3_n8), 
        .Z(prince_rounds_mul_input_s3[11]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_12_U1 ( .A(
        prince_rounds_sub_Result_s3[12]), .B(
        prince_rounds_SR_Inv_Result_s3[12]), .S(prince_rounds_S_Sinv_mul3_n8), 
        .Z(prince_rounds_mul_input_s3[12]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_13_U1 ( .A(
        prince_rounds_sub_Result_s3[13]), .B(
        prince_rounds_SR_Inv_Result_s3[13]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[13]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_14_U1 ( .A(
        prince_rounds_sub_Result_s3[14]), .B(
        prince_rounds_SR_Inv_Result_s3[14]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[14]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_15_U1 ( .A(
        prince_rounds_sub_Result_s3[15]), .B(
        prince_rounds_SR_Inv_Result_s3[15]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[15]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_16_U1 ( .A(
        prince_rounds_sub_Result_s3[16]), .B(
        prince_rounds_SR_Inv_Result_s3[16]), .S(prince_rounds_S_Sinv_mul3_n8), 
        .Z(prince_rounds_mul_input_s3[16]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_17_U1 ( .A(
        prince_rounds_sub_Result_s3[17]), .B(
        prince_rounds_SR_Inv_Result_s3[17]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[17]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_18_U1 ( .A(
        prince_rounds_sub_Result_s3[18]), .B(
        prince_rounds_SR_Inv_Result_s3[18]), .S(prince_rounds_S_Sinv_mul3_n8), 
        .Z(prince_rounds_mul_input_s3[18]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_19_U1 ( .A(
        prince_rounds_sub_Result_s3[19]), .B(
        prince_rounds_SR_Inv_Result_s3[19]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[19]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_20_U1 ( .A(
        prince_rounds_sub_Result_s3[20]), .B(
        prince_rounds_SR_Inv_Result_s3[20]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[20]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_21_U1 ( .A(
        prince_rounds_sub_Result_s3[21]), .B(
        prince_rounds_SR_Inv_Result_s3[21]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[21]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_22_U1 ( .A(
        prince_rounds_sub_Result_s3[22]), .B(
        prince_rounds_SR_Inv_Result_s3[22]), .S(prince_rounds_S_Sinv_mul3_n8), 
        .Z(prince_rounds_mul_input_s3[22]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_23_U1 ( .A(
        prince_rounds_sub_Result_s3[23]), .B(
        prince_rounds_SR_Inv_Result_s3[23]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[23]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_24_U1 ( .A(
        prince_rounds_sub_Result_s3[24]), .B(
        prince_rounds_SR_Inv_Result_s3[24]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[24]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_25_U1 ( .A(
        prince_rounds_sub_Result_s3[25]), .B(
        prince_rounds_SR_Inv_Result_s3[25]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[25]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_26_U1 ( .A(
        prince_rounds_sub_Result_s3[26]), .B(
        prince_rounds_SR_Inv_Result_s3[26]), .S(prince_rounds_S_Sinv_mul3_n8), 
        .Z(prince_rounds_mul_input_s3[26]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_27_U1 ( .A(
        prince_rounds_sub_Result_s3[27]), .B(
        prince_rounds_SR_Inv_Result_s3[27]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[27]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_28_U1 ( .A(
        prince_rounds_sub_Result_s3[28]), .B(
        prince_rounds_SR_Inv_Result_s3[28]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[28]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_29_U1 ( .A(
        prince_rounds_sub_Result_s3[29]), .B(
        prince_rounds_SR_Inv_Result_s3[29]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[29]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_30_U1 ( .A(
        prince_rounds_sub_Result_s3[30]), .B(
        prince_rounds_SR_Inv_Result_s3[30]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[30]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_31_U1 ( .A(
        prince_rounds_sub_Result_s3[31]), .B(
        prince_rounds_SR_Inv_Result_s3[31]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[31]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_32_U1 ( .A(
        prince_rounds_sub_Result_s3[32]), .B(
        prince_rounds_SR_Inv_Result_s3[32]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[32]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_33_U1 ( .A(
        prince_rounds_sub_Result_s3[33]), .B(
        prince_rounds_SR_Inv_Result_s3[33]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[33]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_34_U1 ( .A(
        prince_rounds_sub_Result_s3[34]), .B(
        prince_rounds_SR_Inv_Result_s3[34]), .S(prince_rounds_S_Sinv_mul3_n8), 
        .Z(prince_rounds_mul_input_s3[34]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_35_U1 ( .A(
        prince_rounds_sub_Result_s3[35]), .B(
        prince_rounds_SR_Inv_Result_s3[35]), .S(prince_rounds_S_Sinv_mul3_n6), 
        .Z(prince_rounds_mul_input_s3[35]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_36_U1 ( .A(
        prince_rounds_sub_Result_s3[36]), .B(
        prince_rounds_SR_Inv_Result_s3[36]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s3[36]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_37_U1 ( .A(
        prince_rounds_sub_Result_s3[37]), .B(
        prince_rounds_SR_Inv_Result_s3[37]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s3[37]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_38_U1 ( .A(
        prince_rounds_sub_Result_s3[38]), .B(
        prince_rounds_SR_Inv_Result_s3[38]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s3[38]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_39_U1 ( .A(
        prince_rounds_sub_Result_s3[39]), .B(
        prince_rounds_SR_Inv_Result_s3[39]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s3[39]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_40_U1 ( .A(
        prince_rounds_sub_Result_s3[40]), .B(
        prince_rounds_SR_Inv_Result_s3[40]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s3[40]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_41_U1 ( .A(
        prince_rounds_sub_Result_s3[41]), .B(
        prince_rounds_SR_Inv_Result_s3[41]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s3[41]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_42_U1 ( .A(
        prince_rounds_sub_Result_s3[42]), .B(
        prince_rounds_SR_Inv_Result_s3[42]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s3[42]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_43_U1 ( .A(
        prince_rounds_sub_Result_s3[43]), .B(
        prince_rounds_SR_Inv_Result_s3[43]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s3[43]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_44_U1 ( .A(
        prince_rounds_sub_Result_s3[44]), .B(
        prince_rounds_SR_Inv_Result_s3[44]), .S(prince_rounds_S_Sinv_mul3_n7), 
        .Z(prince_rounds_mul_input_s3[44]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_45_U1 ( .A(
        prince_rounds_sub_Result_s3[45]), .B(
        prince_rounds_SR_Inv_Result_s3[45]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s3[45]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_46_U1 ( .A(
        prince_rounds_sub_Result_s3[46]), .B(
        prince_rounds_SR_Inv_Result_s3[46]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s3[46]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_47_U1 ( .A(
        prince_rounds_sub_Result_s3[47]), .B(
        prince_rounds_SR_Inv_Result_s3[47]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s3[47]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_48_U1 ( .A(
        prince_rounds_sub_Result_s3[48]), .B(
        prince_rounds_SR_Inv_Result_s3[48]), .S(prince_rounds_S_Sinv_mul3_n7), 
        .Z(prince_rounds_mul_input_s3[48]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_49_U1 ( .A(
        prince_rounds_sub_Result_s3[49]), .B(
        prince_rounds_SR_Inv_Result_s3[49]), .S(prince_rounds_S_Sinv_mul3_n7), 
        .Z(prince_rounds_mul_input_s3[49]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_50_U1 ( .A(
        prince_rounds_sub_Result_s3[50]), .B(
        prince_rounds_SR_Inv_Result_s3[50]), .S(prince_rounds_S_Sinv_mul3_n7), 
        .Z(prince_rounds_mul_input_s3[50]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_51_U1 ( .A(
        prince_rounds_sub_Result_s3[51]), .B(
        prince_rounds_SR_Inv_Result_s3[51]), .S(prince_rounds_S_Sinv_mul3_n7), 
        .Z(prince_rounds_mul_input_s3[51]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_52_U1 ( .A(
        prince_rounds_sub_Result_s3[52]), .B(
        prince_rounds_SR_Inv_Result_s3[52]), .S(prince_rounds_S_Sinv_mul3_n7), 
        .Z(prince_rounds_mul_input_s3[52]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_53_U1 ( .A(
        prince_rounds_sub_Result_s3[53]), .B(
        prince_rounds_SR_Inv_Result_s3[53]), .S(prince_rounds_S_Sinv_mul3_n7), 
        .Z(prince_rounds_mul_input_s3[53]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_54_U1 ( .A(
        prince_rounds_sub_Result_s3[54]), .B(
        prince_rounds_SR_Inv_Result_s3[54]), .S(prince_rounds_S_Sinv_mul3_n7), 
        .Z(prince_rounds_mul_input_s3[54]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_55_U1 ( .A(
        prince_rounds_sub_Result_s3[55]), .B(
        prince_rounds_SR_Inv_Result_s3[55]), .S(prince_rounds_S_Sinv_mul3_n7), 
        .Z(prince_rounds_mul_input_s3[55]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_56_U1 ( .A(
        prince_rounds_sub_Result_s3[56]), .B(
        prince_rounds_SR_Inv_Result_s3[56]), .S(prince_rounds_S_Sinv_mul3_n7), 
        .Z(prince_rounds_mul_input_s3[56]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_57_U1 ( .A(
        prince_rounds_sub_Result_s3[57]), .B(
        prince_rounds_SR_Inv_Result_s3[57]), .S(prince_rounds_S_Sinv_mul3_n7), 
        .Z(prince_rounds_mul_input_s3[57]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_58_U1 ( .A(
        prince_rounds_sub_Result_s3[58]), .B(
        prince_rounds_SR_Inv_Result_s3[58]), .S(prince_rounds_S_Sinv_mul3_n7), 
        .Z(prince_rounds_mul_input_s3[58]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_59_U1 ( .A(
        prince_rounds_sub_Result_s3[59]), .B(
        prince_rounds_SR_Inv_Result_s3[59]), .S(prince_rounds_S_Sinv_mul3_n7), 
        .Z(prince_rounds_mul_input_s3[59]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_60_U1 ( .A(
        prince_rounds_sub_Result_s3[60]), .B(
        prince_rounds_SR_Inv_Result_s3[60]), .S(prince_rounds_S_Sinv_mul3_n7), 
        .Z(prince_rounds_mul_input_s3[60]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_61_U1 ( .A(
        prince_rounds_sub_Result_s3[61]), .B(
        prince_rounds_SR_Inv_Result_s3[61]), .S(prince_rounds_S_Sinv_mul3_n7), 
        .Z(prince_rounds_mul_input_s3[61]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_62_U1 ( .A(
        prince_rounds_sub_Result_s3[62]), .B(
        prince_rounds_SR_Inv_Result_s3[62]), .S(prince_rounds_S_Sinv_mul3_n7), 
        .Z(prince_rounds_mul_input_s3[62]) );
  MUX2_X1 prince_rounds_S_Sinv_mul3_MUXInst_63_U1 ( .A(
        prince_rounds_sub_Result_s3[63]), .B(
        prince_rounds_SR_Inv_Result_s3[63]), .S(roundEnd_Select_Signal), .Z(
        prince_rounds_mul_input_s3[63]) );
  XNOR2_X1 prince_rounds_mul_s1_U96 ( .A(prince_rounds_mul_input_s1[13]), .B(
        prince_rounds_mul_s1_n96), .ZN(prince_rounds_mul_result_s1[9]) );
  XNOR2_X1 prince_rounds_mul_s1_U95 ( .A(prince_rounds_mul_input_s1[0]), .B(
        prince_rounds_mul_s1_n95), .ZN(prince_rounds_mul_result_s1[8]) );
  XNOR2_X1 prince_rounds_mul_s1_U94 ( .A(prince_rounds_mul_input_s1[11]), .B(
        prince_rounds_mul_s1_n94), .ZN(prince_rounds_mul_result_s1[7]) );
  XNOR2_X1 prince_rounds_mul_s1_U93 ( .A(prince_rounds_mul_input_s1[10]), .B(
        prince_rounds_mul_s1_n93), .ZN(prince_rounds_mul_result_s1[6]) );
  XNOR2_X1 prince_rounds_mul_s1_U92 ( .A(prince_rounds_mul_input_s1[51]), .B(
        prince_rounds_mul_s1_n92), .ZN(prince_rounds_mul_result_s1[63]) );
  XNOR2_X1 prince_rounds_mul_s1_U91 ( .A(prince_rounds_mul_input_s1[50]), .B(
        prince_rounds_mul_s1_n91), .ZN(prince_rounds_mul_result_s1[62]) );
  XNOR2_X1 prince_rounds_mul_s1_U90 ( .A(prince_rounds_mul_input_s1[49]), .B(
        prince_rounds_mul_s1_n90), .ZN(prince_rounds_mul_result_s1[61]) );
  XNOR2_X1 prince_rounds_mul_s1_U89 ( .A(prince_rounds_mul_input_s1[52]), .B(
        prince_rounds_mul_s1_n89), .ZN(prince_rounds_mul_result_s1[60]) );
  XNOR2_X1 prince_rounds_mul_s1_U88 ( .A(prince_rounds_mul_input_s1[9]), .B(
        prince_rounds_mul_s1_n96), .ZN(prince_rounds_mul_result_s1[5]) );
  XNOR2_X1 prince_rounds_mul_s1_U87 ( .A(prince_rounds_mul_input_s1[1]), .B(
        prince_rounds_mul_input_s1[5]), .ZN(prince_rounds_mul_s1_n96) );
  XNOR2_X1 prince_rounds_mul_s1_U86 ( .A(prince_rounds_mul_input_s1[63]), .B(
        prince_rounds_mul_s1_n92), .ZN(prince_rounds_mul_result_s1[59]) );
  XNOR2_X1 prince_rounds_mul_s1_U85 ( .A(prince_rounds_mul_input_s1[55]), .B(
        prince_rounds_mul_input_s1[59]), .ZN(prince_rounds_mul_s1_n92) );
  XNOR2_X1 prince_rounds_mul_s1_U84 ( .A(prince_rounds_mul_input_s1[54]), .B(
        prince_rounds_mul_s1_n88), .ZN(prince_rounds_mul_result_s1[58]) );
  XNOR2_X1 prince_rounds_mul_s1_U83 ( .A(prince_rounds_mul_input_s1[61]), .B(
        prince_rounds_mul_s1_n87), .ZN(prince_rounds_mul_result_s1[57]) );
  XNOR2_X1 prince_rounds_mul_s1_U82 ( .A(prince_rounds_mul_input_s1[48]), .B(
        prince_rounds_mul_s1_n89), .ZN(prince_rounds_mul_result_s1[56]) );
  XNOR2_X1 prince_rounds_mul_s1_U81 ( .A(prince_rounds_mul_input_s1[56]), .B(
        prince_rounds_mul_input_s1[60]), .ZN(prince_rounds_mul_s1_n89) );
  XNOR2_X1 prince_rounds_mul_s1_U80 ( .A(prince_rounds_mul_input_s1[59]), .B(
        prince_rounds_mul_s1_n86), .ZN(prince_rounds_mul_result_s1[55]) );
  XNOR2_X1 prince_rounds_mul_s1_U79 ( .A(prince_rounds_mul_input_s1[58]), .B(
        prince_rounds_mul_s1_n91), .ZN(prince_rounds_mul_result_s1[54]) );
  XNOR2_X1 prince_rounds_mul_s1_U78 ( .A(prince_rounds_mul_input_s1[62]), .B(
        prince_rounds_mul_input_s1[54]), .ZN(prince_rounds_mul_s1_n91) );
  XNOR2_X1 prince_rounds_mul_s1_U77 ( .A(prince_rounds_mul_input_s1[57]), .B(
        prince_rounds_mul_s1_n87), .ZN(prince_rounds_mul_result_s1[53]) );
  XNOR2_X1 prince_rounds_mul_s1_U76 ( .A(prince_rounds_mul_input_s1[53]), .B(
        prince_rounds_mul_input_s1[49]), .ZN(prince_rounds_mul_s1_n87) );
  XNOR2_X1 prince_rounds_mul_s1_U75 ( .A(prince_rounds_mul_input_s1[60]), .B(
        prince_rounds_mul_s1_n85), .ZN(prince_rounds_mul_result_s1[52]) );
  XNOR2_X1 prince_rounds_mul_s1_U74 ( .A(prince_rounds_mul_input_s1[55]), .B(
        prince_rounds_mul_s1_n86), .ZN(prince_rounds_mul_result_s1[51]) );
  XNOR2_X1 prince_rounds_mul_s1_U73 ( .A(prince_rounds_mul_input_s1[51]), .B(
        prince_rounds_mul_input_s1[63]), .ZN(prince_rounds_mul_s1_n86) );
  XNOR2_X1 prince_rounds_mul_s1_U72 ( .A(prince_rounds_mul_input_s1[62]), .B(
        prince_rounds_mul_s1_n88), .ZN(prince_rounds_mul_result_s1[50]) );
  XNOR2_X1 prince_rounds_mul_s1_U71 ( .A(prince_rounds_mul_input_s1[50]), .B(
        prince_rounds_mul_input_s1[58]), .ZN(prince_rounds_mul_s1_n88) );
  XNOR2_X1 prince_rounds_mul_s1_U70 ( .A(prince_rounds_mul_input_s1[12]), .B(
        prince_rounds_mul_s1_n84), .ZN(prince_rounds_mul_result_s1[4]) );
  XNOR2_X1 prince_rounds_mul_s1_U69 ( .A(prince_rounds_mul_input_s1[53]), .B(
        prince_rounds_mul_s1_n90), .ZN(prince_rounds_mul_result_s1[49]) );
  XNOR2_X1 prince_rounds_mul_s1_U68 ( .A(prince_rounds_mul_input_s1[57]), .B(
        prince_rounds_mul_input_s1[61]), .ZN(prince_rounds_mul_s1_n90) );
  XNOR2_X1 prince_rounds_mul_s1_U67 ( .A(prince_rounds_mul_input_s1[56]), .B(
        prince_rounds_mul_s1_n85), .ZN(prince_rounds_mul_result_s1[48]) );
  XNOR2_X1 prince_rounds_mul_s1_U66 ( .A(prince_rounds_mul_input_s1[52]), .B(
        prince_rounds_mul_input_s1[48]), .ZN(prince_rounds_mul_s1_n85) );
  XNOR2_X1 prince_rounds_mul_s1_U65 ( .A(prince_rounds_mul_input_s1[39]), .B(
        prince_rounds_mul_s1_n83), .ZN(prince_rounds_mul_result_s1[47]) );
  XNOR2_X1 prince_rounds_mul_s1_U64 ( .A(prince_rounds_mul_input_s1[34]), .B(
        prince_rounds_mul_s1_n82), .ZN(prince_rounds_mul_result_s1[46]) );
  XNOR2_X1 prince_rounds_mul_s1_U63 ( .A(prince_rounds_mul_input_s1[33]), .B(
        prince_rounds_mul_s1_n81), .ZN(prince_rounds_mul_result_s1[45]) );
  XNOR2_X1 prince_rounds_mul_s1_U62 ( .A(prince_rounds_mul_input_s1[32]), .B(
        prince_rounds_mul_s1_n80), .ZN(prince_rounds_mul_result_s1[44]) );
  XNOR2_X1 prince_rounds_mul_s1_U61 ( .A(prince_rounds_mul_input_s1[35]), .B(
        prince_rounds_mul_s1_n83), .ZN(prince_rounds_mul_result_s1[43]) );
  XNOR2_X1 prince_rounds_mul_s1_U60 ( .A(prince_rounds_mul_input_s1[43]), .B(
        prince_rounds_mul_input_s1[47]), .ZN(prince_rounds_mul_s1_n83) );
  XNOR2_X1 prince_rounds_mul_s1_U59 ( .A(prince_rounds_mul_input_s1[46]), .B(
        prince_rounds_mul_s1_n82), .ZN(prince_rounds_mul_result_s1[42]) );
  XNOR2_X1 prince_rounds_mul_s1_U58 ( .A(prince_rounds_mul_input_s1[38]), .B(
        prince_rounds_mul_input_s1[42]), .ZN(prince_rounds_mul_s1_n82) );
  XNOR2_X1 prince_rounds_mul_s1_U57 ( .A(prince_rounds_mul_input_s1[37]), .B(
        prince_rounds_mul_s1_n79), .ZN(prince_rounds_mul_result_s1[41]) );
  XNOR2_X1 prince_rounds_mul_s1_U56 ( .A(prince_rounds_mul_input_s1[44]), .B(
        prince_rounds_mul_s1_n78), .ZN(prince_rounds_mul_result_s1[40]) );
  XNOR2_X1 prince_rounds_mul_s1_U55 ( .A(prince_rounds_mul_input_s1[7]), .B(
        prince_rounds_mul_s1_n94), .ZN(prince_rounds_mul_result_s1[3]) );
  XNOR2_X1 prince_rounds_mul_s1_U54 ( .A(prince_rounds_mul_input_s1[15]), .B(
        prince_rounds_mul_input_s1[3]), .ZN(prince_rounds_mul_s1_n94) );
  XNOR2_X1 prince_rounds_mul_s1_U53 ( .A(prince_rounds_mul_input_s1[47]), .B(
        prince_rounds_mul_s1_n77), .ZN(prince_rounds_mul_result_s1[39]) );
  XNOR2_X1 prince_rounds_mul_s1_U52 ( .A(prince_rounds_mul_input_s1[42]), .B(
        prince_rounds_mul_s1_n76), .ZN(prince_rounds_mul_result_s1[38]) );
  XNOR2_X1 prince_rounds_mul_s1_U51 ( .A(prince_rounds_mul_input_s1[41]), .B(
        prince_rounds_mul_s1_n81), .ZN(prince_rounds_mul_result_s1[37]) );
  XNOR2_X1 prince_rounds_mul_s1_U50 ( .A(prince_rounds_mul_input_s1[45]), .B(
        prince_rounds_mul_input_s1[37]), .ZN(prince_rounds_mul_s1_n81) );
  XNOR2_X1 prince_rounds_mul_s1_U49 ( .A(prince_rounds_mul_input_s1[40]), .B(
        prince_rounds_mul_s1_n78), .ZN(prince_rounds_mul_result_s1[36]) );
  XNOR2_X1 prince_rounds_mul_s1_U48 ( .A(prince_rounds_mul_input_s1[36]), .B(
        prince_rounds_mul_input_s1[32]), .ZN(prince_rounds_mul_s1_n78) );
  XNOR2_X1 prince_rounds_mul_s1_U47 ( .A(prince_rounds_mul_input_s1[43]), .B(
        prince_rounds_mul_s1_n77), .ZN(prince_rounds_mul_result_s1[35]) );
  XNOR2_X1 prince_rounds_mul_s1_U46 ( .A(prince_rounds_mul_input_s1[39]), .B(
        prince_rounds_mul_input_s1[35]), .ZN(prince_rounds_mul_s1_n77) );
  XNOR2_X1 prince_rounds_mul_s1_U45 ( .A(prince_rounds_mul_input_s1[38]), .B(
        prince_rounds_mul_s1_n76), .ZN(prince_rounds_mul_result_s1[34]) );
  XNOR2_X1 prince_rounds_mul_s1_U44 ( .A(prince_rounds_mul_input_s1[34]), .B(
        prince_rounds_mul_input_s1[46]), .ZN(prince_rounds_mul_s1_n76) );
  XNOR2_X1 prince_rounds_mul_s1_U43 ( .A(prince_rounds_mul_input_s1[45]), .B(
        prince_rounds_mul_s1_n79), .ZN(prince_rounds_mul_result_s1[33]) );
  XNOR2_X1 prince_rounds_mul_s1_U42 ( .A(prince_rounds_mul_input_s1[33]), .B(
        prince_rounds_mul_input_s1[41]), .ZN(prince_rounds_mul_s1_n79) );
  XNOR2_X1 prince_rounds_mul_s1_U41 ( .A(prince_rounds_mul_input_s1[36]), .B(
        prince_rounds_mul_s1_n80), .ZN(prince_rounds_mul_result_s1[32]) );
  XNOR2_X1 prince_rounds_mul_s1_U40 ( .A(prince_rounds_mul_input_s1[40]), .B(
        prince_rounds_mul_input_s1[44]), .ZN(prince_rounds_mul_s1_n80) );
  XNOR2_X1 prince_rounds_mul_s1_U39 ( .A(prince_rounds_mul_input_s1[23]), .B(
        prince_rounds_mul_s1_n75), .ZN(prince_rounds_mul_result_s1[31]) );
  XNOR2_X1 prince_rounds_mul_s1_U38 ( .A(prince_rounds_mul_input_s1[18]), .B(
        prince_rounds_mul_s1_n74), .ZN(prince_rounds_mul_result_s1[30]) );
  XNOR2_X1 prince_rounds_mul_s1_U37 ( .A(prince_rounds_mul_input_s1[14]), .B(
        prince_rounds_mul_s1_n73), .ZN(prince_rounds_mul_result_s1[2]) );
  XNOR2_X1 prince_rounds_mul_s1_U36 ( .A(prince_rounds_mul_input_s1[17]), .B(
        prince_rounds_mul_s1_n72), .ZN(prince_rounds_mul_result_s1[29]) );
  XNOR2_X1 prince_rounds_mul_s1_U35 ( .A(prince_rounds_mul_input_s1[16]), .B(
        prince_rounds_mul_s1_n71), .ZN(prince_rounds_mul_result_s1[28]) );
  XNOR2_X1 prince_rounds_mul_s1_U34 ( .A(prince_rounds_mul_input_s1[19]), .B(
        prince_rounds_mul_s1_n75), .ZN(prince_rounds_mul_result_s1[27]) );
  XNOR2_X1 prince_rounds_mul_s1_U33 ( .A(prince_rounds_mul_input_s1[27]), .B(
        prince_rounds_mul_input_s1[31]), .ZN(prince_rounds_mul_s1_n75) );
  XNOR2_X1 prince_rounds_mul_s1_U32 ( .A(prince_rounds_mul_input_s1[30]), .B(
        prince_rounds_mul_s1_n74), .ZN(prince_rounds_mul_result_s1[26]) );
  XNOR2_X1 prince_rounds_mul_s1_U31 ( .A(prince_rounds_mul_input_s1[22]), .B(
        prince_rounds_mul_input_s1[26]), .ZN(prince_rounds_mul_s1_n74) );
  XNOR2_X1 prince_rounds_mul_s1_U30 ( .A(prince_rounds_mul_input_s1[21]), .B(
        prince_rounds_mul_s1_n70), .ZN(prince_rounds_mul_result_s1[25]) );
  XNOR2_X1 prince_rounds_mul_s1_U29 ( .A(prince_rounds_mul_input_s1[28]), .B(
        prince_rounds_mul_s1_n69), .ZN(prince_rounds_mul_result_s1[24]) );
  XNOR2_X1 prince_rounds_mul_s1_U28 ( .A(prince_rounds_mul_input_s1[31]), .B(
        prince_rounds_mul_s1_n68), .ZN(prince_rounds_mul_result_s1[23]) );
  XNOR2_X1 prince_rounds_mul_s1_U27 ( .A(prince_rounds_mul_input_s1[26]), .B(
        prince_rounds_mul_s1_n67), .ZN(prince_rounds_mul_result_s1[22]) );
  XNOR2_X1 prince_rounds_mul_s1_U26 ( .A(prince_rounds_mul_input_s1[25]), .B(
        prince_rounds_mul_s1_n72), .ZN(prince_rounds_mul_result_s1[21]) );
  XNOR2_X1 prince_rounds_mul_s1_U25 ( .A(prince_rounds_mul_input_s1[29]), .B(
        prince_rounds_mul_input_s1[21]), .ZN(prince_rounds_mul_s1_n72) );
  XNOR2_X1 prince_rounds_mul_s1_U24 ( .A(prince_rounds_mul_input_s1[24]), .B(
        prince_rounds_mul_s1_n69), .ZN(prince_rounds_mul_result_s1[20]) );
  XNOR2_X1 prince_rounds_mul_s1_U23 ( .A(prince_rounds_mul_input_s1[20]), .B(
        prince_rounds_mul_input_s1[16]), .ZN(prince_rounds_mul_s1_n69) );
  XNOR2_X1 prince_rounds_mul_s1_U22 ( .A(prince_rounds_mul_input_s1[5]), .B(
        prince_rounds_mul_s1_n66), .ZN(prince_rounds_mul_result_s1[1]) );
  XNOR2_X1 prince_rounds_mul_s1_U21 ( .A(prince_rounds_mul_input_s1[27]), .B(
        prince_rounds_mul_s1_n68), .ZN(prince_rounds_mul_result_s1[19]) );
  XNOR2_X1 prince_rounds_mul_s1_U20 ( .A(prince_rounds_mul_input_s1[23]), .B(
        prince_rounds_mul_input_s1[19]), .ZN(prince_rounds_mul_s1_n68) );
  XNOR2_X1 prince_rounds_mul_s1_U19 ( .A(prince_rounds_mul_input_s1[22]), .B(
        prince_rounds_mul_s1_n67), .ZN(prince_rounds_mul_result_s1[18]) );
  XNOR2_X1 prince_rounds_mul_s1_U18 ( .A(prince_rounds_mul_input_s1[18]), .B(
        prince_rounds_mul_input_s1[30]), .ZN(prince_rounds_mul_s1_n67) );
  XNOR2_X1 prince_rounds_mul_s1_U17 ( .A(prince_rounds_mul_input_s1[29]), .B(
        prince_rounds_mul_s1_n70), .ZN(prince_rounds_mul_result_s1[17]) );
  XNOR2_X1 prince_rounds_mul_s1_U16 ( .A(prince_rounds_mul_input_s1[17]), .B(
        prince_rounds_mul_input_s1[25]), .ZN(prince_rounds_mul_s1_n70) );
  XNOR2_X1 prince_rounds_mul_s1_U15 ( .A(prince_rounds_mul_input_s1[20]), .B(
        prince_rounds_mul_s1_n71), .ZN(prince_rounds_mul_result_s1[16]) );
  XNOR2_X1 prince_rounds_mul_s1_U14 ( .A(prince_rounds_mul_input_s1[24]), .B(
        prince_rounds_mul_input_s1[28]), .ZN(prince_rounds_mul_s1_n71) );
  XNOR2_X1 prince_rounds_mul_s1_U13 ( .A(prince_rounds_mul_input_s1[3]), .B(
        prince_rounds_mul_s1_n65), .ZN(prince_rounds_mul_result_s1[15]) );
  XNOR2_X1 prince_rounds_mul_s1_U12 ( .A(prince_rounds_mul_input_s1[2]), .B(
        prince_rounds_mul_s1_n93), .ZN(prince_rounds_mul_result_s1[14]) );
  XNOR2_X1 prince_rounds_mul_s1_U11 ( .A(prince_rounds_mul_input_s1[6]), .B(
        prince_rounds_mul_input_s1[14]), .ZN(prince_rounds_mul_s1_n93) );
  XNOR2_X1 prince_rounds_mul_s1_U10 ( .A(prince_rounds_mul_input_s1[1]), .B(
        prince_rounds_mul_s1_n66), .ZN(prince_rounds_mul_result_s1[13]) );
  XNOR2_X1 prince_rounds_mul_s1_U9 ( .A(prince_rounds_mul_input_s1[13]), .B(
        prince_rounds_mul_input_s1[9]), .ZN(prince_rounds_mul_s1_n66) );
  XNOR2_X1 prince_rounds_mul_s1_U8 ( .A(prince_rounds_mul_input_s1[4]), .B(
        prince_rounds_mul_s1_n95), .ZN(prince_rounds_mul_result_s1[12]) );
  XNOR2_X1 prince_rounds_mul_s1_U7 ( .A(prince_rounds_mul_input_s1[8]), .B(
        prince_rounds_mul_input_s1[12]), .ZN(prince_rounds_mul_s1_n95) );
  XNOR2_X1 prince_rounds_mul_s1_U6 ( .A(prince_rounds_mul_input_s1[15]), .B(
        prince_rounds_mul_s1_n65), .ZN(prince_rounds_mul_result_s1[11]) );
  XNOR2_X1 prince_rounds_mul_s1_U5 ( .A(prince_rounds_mul_input_s1[11]), .B(
        prince_rounds_mul_input_s1[7]), .ZN(prince_rounds_mul_s1_n65) );
  XNOR2_X1 prince_rounds_mul_s1_U4 ( .A(prince_rounds_mul_input_s1[6]), .B(
        prince_rounds_mul_s1_n73), .ZN(prince_rounds_mul_result_s1[10]) );
  XNOR2_X1 prince_rounds_mul_s1_U3 ( .A(prince_rounds_mul_input_s1[10]), .B(
        prince_rounds_mul_input_s1[2]), .ZN(prince_rounds_mul_s1_n73) );
  XNOR2_X1 prince_rounds_mul_s1_U2 ( .A(prince_rounds_mul_input_s1[8]), .B(
        prince_rounds_mul_s1_n84), .ZN(prince_rounds_mul_result_s1[0]) );
  XNOR2_X1 prince_rounds_mul_s1_U1 ( .A(prince_rounds_mul_input_s1[0]), .B(
        prince_rounds_mul_input_s1[4]), .ZN(prince_rounds_mul_s1_n84) );
  XNOR2_X1 prince_rounds_mul_s2_U96 ( .A(prince_rounds_mul_input_s2[13]), .B(
        prince_rounds_mul_s2_n96), .ZN(prince_rounds_mul_result_s2[9]) );
  XNOR2_X1 prince_rounds_mul_s2_U95 ( .A(prince_rounds_mul_input_s2[0]), .B(
        prince_rounds_mul_s2_n95), .ZN(prince_rounds_mul_result_s2[8]) );
  XNOR2_X1 prince_rounds_mul_s2_U94 ( .A(prince_rounds_mul_input_s2[11]), .B(
        prince_rounds_mul_s2_n94), .ZN(prince_rounds_mul_result_s2[7]) );
  XNOR2_X1 prince_rounds_mul_s2_U93 ( .A(prince_rounds_mul_input_s2[10]), .B(
        prince_rounds_mul_s2_n93), .ZN(prince_rounds_mul_result_s2[6]) );
  XNOR2_X1 prince_rounds_mul_s2_U92 ( .A(prince_rounds_mul_input_s2[51]), .B(
        prince_rounds_mul_s2_n92), .ZN(prince_rounds_mul_result_s2[63]) );
  XNOR2_X1 prince_rounds_mul_s2_U91 ( .A(prince_rounds_mul_input_s2[50]), .B(
        prince_rounds_mul_s2_n91), .ZN(prince_rounds_mul_result_s2[62]) );
  XNOR2_X1 prince_rounds_mul_s2_U90 ( .A(prince_rounds_mul_input_s2[49]), .B(
        prince_rounds_mul_s2_n90), .ZN(prince_rounds_mul_result_s2[61]) );
  XNOR2_X1 prince_rounds_mul_s2_U89 ( .A(prince_rounds_mul_input_s2[52]), .B(
        prince_rounds_mul_s2_n89), .ZN(prince_rounds_mul_result_s2[60]) );
  XNOR2_X1 prince_rounds_mul_s2_U88 ( .A(prince_rounds_mul_input_s2[9]), .B(
        prince_rounds_mul_s2_n96), .ZN(prince_rounds_mul_result_s2[5]) );
  XNOR2_X1 prince_rounds_mul_s2_U87 ( .A(prince_rounds_mul_input_s2[1]), .B(
        prince_rounds_mul_input_s2[5]), .ZN(prince_rounds_mul_s2_n96) );
  XNOR2_X1 prince_rounds_mul_s2_U86 ( .A(prince_rounds_mul_input_s2[63]), .B(
        prince_rounds_mul_s2_n92), .ZN(prince_rounds_mul_result_s2[59]) );
  XNOR2_X1 prince_rounds_mul_s2_U85 ( .A(prince_rounds_mul_input_s2[55]), .B(
        prince_rounds_mul_input_s2[59]), .ZN(prince_rounds_mul_s2_n92) );
  XNOR2_X1 prince_rounds_mul_s2_U84 ( .A(prince_rounds_mul_input_s2[54]), .B(
        prince_rounds_mul_s2_n88), .ZN(prince_rounds_mul_result_s2[58]) );
  XNOR2_X1 prince_rounds_mul_s2_U83 ( .A(prince_rounds_mul_input_s2[61]), .B(
        prince_rounds_mul_s2_n87), .ZN(prince_rounds_mul_result_s2[57]) );
  XNOR2_X1 prince_rounds_mul_s2_U82 ( .A(prince_rounds_mul_input_s2[48]), .B(
        prince_rounds_mul_s2_n89), .ZN(prince_rounds_mul_result_s2[56]) );
  XNOR2_X1 prince_rounds_mul_s2_U81 ( .A(prince_rounds_mul_input_s2[56]), .B(
        prince_rounds_mul_input_s2[60]), .ZN(prince_rounds_mul_s2_n89) );
  XNOR2_X1 prince_rounds_mul_s2_U80 ( .A(prince_rounds_mul_input_s2[59]), .B(
        prince_rounds_mul_s2_n86), .ZN(prince_rounds_mul_result_s2[55]) );
  XNOR2_X1 prince_rounds_mul_s2_U79 ( .A(prince_rounds_mul_input_s2[58]), .B(
        prince_rounds_mul_s2_n91), .ZN(prince_rounds_mul_result_s2[54]) );
  XNOR2_X1 prince_rounds_mul_s2_U78 ( .A(prince_rounds_mul_input_s2[62]), .B(
        prince_rounds_mul_input_s2[54]), .ZN(prince_rounds_mul_s2_n91) );
  XNOR2_X1 prince_rounds_mul_s2_U77 ( .A(prince_rounds_mul_input_s2[57]), .B(
        prince_rounds_mul_s2_n87), .ZN(prince_rounds_mul_result_s2[53]) );
  XNOR2_X1 prince_rounds_mul_s2_U76 ( .A(prince_rounds_mul_input_s2[53]), .B(
        prince_rounds_mul_input_s2[49]), .ZN(prince_rounds_mul_s2_n87) );
  XNOR2_X1 prince_rounds_mul_s2_U75 ( .A(prince_rounds_mul_input_s2[60]), .B(
        prince_rounds_mul_s2_n85), .ZN(prince_rounds_mul_result_s2[52]) );
  XNOR2_X1 prince_rounds_mul_s2_U74 ( .A(prince_rounds_mul_input_s2[55]), .B(
        prince_rounds_mul_s2_n86), .ZN(prince_rounds_mul_result_s2[51]) );
  XNOR2_X1 prince_rounds_mul_s2_U73 ( .A(prince_rounds_mul_input_s2[51]), .B(
        prince_rounds_mul_input_s2[63]), .ZN(prince_rounds_mul_s2_n86) );
  XNOR2_X1 prince_rounds_mul_s2_U72 ( .A(prince_rounds_mul_input_s2[62]), .B(
        prince_rounds_mul_s2_n88), .ZN(prince_rounds_mul_result_s2[50]) );
  XNOR2_X1 prince_rounds_mul_s2_U71 ( .A(prince_rounds_mul_input_s2[50]), .B(
        prince_rounds_mul_input_s2[58]), .ZN(prince_rounds_mul_s2_n88) );
  XNOR2_X1 prince_rounds_mul_s2_U70 ( .A(prince_rounds_mul_input_s2[12]), .B(
        prince_rounds_mul_s2_n84), .ZN(prince_rounds_mul_result_s2[4]) );
  XNOR2_X1 prince_rounds_mul_s2_U69 ( .A(prince_rounds_mul_input_s2[53]), .B(
        prince_rounds_mul_s2_n90), .ZN(prince_rounds_mul_result_s2[49]) );
  XNOR2_X1 prince_rounds_mul_s2_U68 ( .A(prince_rounds_mul_input_s2[57]), .B(
        prince_rounds_mul_input_s2[61]), .ZN(prince_rounds_mul_s2_n90) );
  XNOR2_X1 prince_rounds_mul_s2_U67 ( .A(prince_rounds_mul_input_s2[56]), .B(
        prince_rounds_mul_s2_n85), .ZN(prince_rounds_mul_result_s2[48]) );
  XNOR2_X1 prince_rounds_mul_s2_U66 ( .A(prince_rounds_mul_input_s2[52]), .B(
        prince_rounds_mul_input_s2[48]), .ZN(prince_rounds_mul_s2_n85) );
  XNOR2_X1 prince_rounds_mul_s2_U65 ( .A(prince_rounds_mul_input_s2[39]), .B(
        prince_rounds_mul_s2_n83), .ZN(prince_rounds_mul_result_s2[47]) );
  XNOR2_X1 prince_rounds_mul_s2_U64 ( .A(prince_rounds_mul_input_s2[34]), .B(
        prince_rounds_mul_s2_n82), .ZN(prince_rounds_mul_result_s2[46]) );
  XNOR2_X1 prince_rounds_mul_s2_U63 ( .A(prince_rounds_mul_input_s2[33]), .B(
        prince_rounds_mul_s2_n81), .ZN(prince_rounds_mul_result_s2[45]) );
  XNOR2_X1 prince_rounds_mul_s2_U62 ( .A(prince_rounds_mul_input_s2[32]), .B(
        prince_rounds_mul_s2_n80), .ZN(prince_rounds_mul_result_s2[44]) );
  XNOR2_X1 prince_rounds_mul_s2_U61 ( .A(prince_rounds_mul_input_s2[35]), .B(
        prince_rounds_mul_s2_n83), .ZN(prince_rounds_mul_result_s2[43]) );
  XNOR2_X1 prince_rounds_mul_s2_U60 ( .A(prince_rounds_mul_input_s2[43]), .B(
        prince_rounds_mul_input_s2[47]), .ZN(prince_rounds_mul_s2_n83) );
  XNOR2_X1 prince_rounds_mul_s2_U59 ( .A(prince_rounds_mul_input_s2[46]), .B(
        prince_rounds_mul_s2_n82), .ZN(prince_rounds_mul_result_s2[42]) );
  XNOR2_X1 prince_rounds_mul_s2_U58 ( .A(prince_rounds_mul_input_s2[38]), .B(
        prince_rounds_mul_input_s2[42]), .ZN(prince_rounds_mul_s2_n82) );
  XNOR2_X1 prince_rounds_mul_s2_U57 ( .A(prince_rounds_mul_input_s2[37]), .B(
        prince_rounds_mul_s2_n79), .ZN(prince_rounds_mul_result_s2[41]) );
  XNOR2_X1 prince_rounds_mul_s2_U56 ( .A(prince_rounds_mul_input_s2[44]), .B(
        prince_rounds_mul_s2_n78), .ZN(prince_rounds_mul_result_s2[40]) );
  XNOR2_X1 prince_rounds_mul_s2_U55 ( .A(prince_rounds_mul_input_s2[7]), .B(
        prince_rounds_mul_s2_n94), .ZN(prince_rounds_mul_result_s2[3]) );
  XNOR2_X1 prince_rounds_mul_s2_U54 ( .A(prince_rounds_mul_input_s2[15]), .B(
        prince_rounds_mul_input_s2[3]), .ZN(prince_rounds_mul_s2_n94) );
  XNOR2_X1 prince_rounds_mul_s2_U53 ( .A(prince_rounds_mul_input_s2[47]), .B(
        prince_rounds_mul_s2_n77), .ZN(prince_rounds_mul_result_s2[39]) );
  XNOR2_X1 prince_rounds_mul_s2_U52 ( .A(prince_rounds_mul_input_s2[42]), .B(
        prince_rounds_mul_s2_n76), .ZN(prince_rounds_mul_result_s2[38]) );
  XNOR2_X1 prince_rounds_mul_s2_U51 ( .A(prince_rounds_mul_input_s2[41]), .B(
        prince_rounds_mul_s2_n81), .ZN(prince_rounds_mul_result_s2[37]) );
  XNOR2_X1 prince_rounds_mul_s2_U50 ( .A(prince_rounds_mul_input_s2[45]), .B(
        prince_rounds_mul_input_s2[37]), .ZN(prince_rounds_mul_s2_n81) );
  XNOR2_X1 prince_rounds_mul_s2_U49 ( .A(prince_rounds_mul_input_s2[40]), .B(
        prince_rounds_mul_s2_n78), .ZN(prince_rounds_mul_result_s2[36]) );
  XNOR2_X1 prince_rounds_mul_s2_U48 ( .A(prince_rounds_mul_input_s2[36]), .B(
        prince_rounds_mul_input_s2[32]), .ZN(prince_rounds_mul_s2_n78) );
  XNOR2_X1 prince_rounds_mul_s2_U47 ( .A(prince_rounds_mul_input_s2[43]), .B(
        prince_rounds_mul_s2_n77), .ZN(prince_rounds_mul_result_s2[35]) );
  XNOR2_X1 prince_rounds_mul_s2_U46 ( .A(prince_rounds_mul_input_s2[39]), .B(
        prince_rounds_mul_input_s2[35]), .ZN(prince_rounds_mul_s2_n77) );
  XNOR2_X1 prince_rounds_mul_s2_U45 ( .A(prince_rounds_mul_input_s2[38]), .B(
        prince_rounds_mul_s2_n76), .ZN(prince_rounds_mul_result_s2[34]) );
  XNOR2_X1 prince_rounds_mul_s2_U44 ( .A(prince_rounds_mul_input_s2[34]), .B(
        prince_rounds_mul_input_s2[46]), .ZN(prince_rounds_mul_s2_n76) );
  XNOR2_X1 prince_rounds_mul_s2_U43 ( .A(prince_rounds_mul_input_s2[45]), .B(
        prince_rounds_mul_s2_n79), .ZN(prince_rounds_mul_result_s2[33]) );
  XNOR2_X1 prince_rounds_mul_s2_U42 ( .A(prince_rounds_mul_input_s2[33]), .B(
        prince_rounds_mul_input_s2[41]), .ZN(prince_rounds_mul_s2_n79) );
  XNOR2_X1 prince_rounds_mul_s2_U41 ( .A(prince_rounds_mul_input_s2[36]), .B(
        prince_rounds_mul_s2_n80), .ZN(prince_rounds_mul_result_s2[32]) );
  XNOR2_X1 prince_rounds_mul_s2_U40 ( .A(prince_rounds_mul_input_s2[40]), .B(
        prince_rounds_mul_input_s2[44]), .ZN(prince_rounds_mul_s2_n80) );
  XNOR2_X1 prince_rounds_mul_s2_U39 ( .A(prince_rounds_mul_input_s2[23]), .B(
        prince_rounds_mul_s2_n75), .ZN(prince_rounds_mul_result_s2[31]) );
  XNOR2_X1 prince_rounds_mul_s2_U38 ( .A(prince_rounds_mul_input_s2[18]), .B(
        prince_rounds_mul_s2_n74), .ZN(prince_rounds_mul_result_s2[30]) );
  XNOR2_X1 prince_rounds_mul_s2_U37 ( .A(prince_rounds_mul_input_s2[14]), .B(
        prince_rounds_mul_s2_n73), .ZN(prince_rounds_mul_result_s2[2]) );
  XNOR2_X1 prince_rounds_mul_s2_U36 ( .A(prince_rounds_mul_input_s2[17]), .B(
        prince_rounds_mul_s2_n72), .ZN(prince_rounds_mul_result_s2[29]) );
  XNOR2_X1 prince_rounds_mul_s2_U35 ( .A(prince_rounds_mul_input_s2[16]), .B(
        prince_rounds_mul_s2_n71), .ZN(prince_rounds_mul_result_s2[28]) );
  XNOR2_X1 prince_rounds_mul_s2_U34 ( .A(prince_rounds_mul_input_s2[19]), .B(
        prince_rounds_mul_s2_n75), .ZN(prince_rounds_mul_result_s2[27]) );
  XNOR2_X1 prince_rounds_mul_s2_U33 ( .A(prince_rounds_mul_input_s2[27]), .B(
        prince_rounds_mul_input_s2[31]), .ZN(prince_rounds_mul_s2_n75) );
  XNOR2_X1 prince_rounds_mul_s2_U32 ( .A(prince_rounds_mul_input_s2[30]), .B(
        prince_rounds_mul_s2_n74), .ZN(prince_rounds_mul_result_s2[26]) );
  XNOR2_X1 prince_rounds_mul_s2_U31 ( .A(prince_rounds_mul_input_s2[22]), .B(
        prince_rounds_mul_input_s2[26]), .ZN(prince_rounds_mul_s2_n74) );
  XNOR2_X1 prince_rounds_mul_s2_U30 ( .A(prince_rounds_mul_input_s2[21]), .B(
        prince_rounds_mul_s2_n70), .ZN(prince_rounds_mul_result_s2[25]) );
  XNOR2_X1 prince_rounds_mul_s2_U29 ( .A(prince_rounds_mul_input_s2[28]), .B(
        prince_rounds_mul_s2_n69), .ZN(prince_rounds_mul_result_s2[24]) );
  XNOR2_X1 prince_rounds_mul_s2_U28 ( .A(prince_rounds_mul_input_s2[31]), .B(
        prince_rounds_mul_s2_n68), .ZN(prince_rounds_mul_result_s2[23]) );
  XNOR2_X1 prince_rounds_mul_s2_U27 ( .A(prince_rounds_mul_input_s2[26]), .B(
        prince_rounds_mul_s2_n67), .ZN(prince_rounds_mul_result_s2[22]) );
  XNOR2_X1 prince_rounds_mul_s2_U26 ( .A(prince_rounds_mul_input_s2[25]), .B(
        prince_rounds_mul_s2_n72), .ZN(prince_rounds_mul_result_s2[21]) );
  XNOR2_X1 prince_rounds_mul_s2_U25 ( .A(prince_rounds_mul_input_s2[29]), .B(
        prince_rounds_mul_input_s2[21]), .ZN(prince_rounds_mul_s2_n72) );
  XNOR2_X1 prince_rounds_mul_s2_U24 ( .A(prince_rounds_mul_input_s2[24]), .B(
        prince_rounds_mul_s2_n69), .ZN(prince_rounds_mul_result_s2[20]) );
  XNOR2_X1 prince_rounds_mul_s2_U23 ( .A(prince_rounds_mul_input_s2[20]), .B(
        prince_rounds_mul_input_s2[16]), .ZN(prince_rounds_mul_s2_n69) );
  XNOR2_X1 prince_rounds_mul_s2_U22 ( .A(prince_rounds_mul_input_s2[5]), .B(
        prince_rounds_mul_s2_n66), .ZN(prince_rounds_mul_result_s2[1]) );
  XNOR2_X1 prince_rounds_mul_s2_U21 ( .A(prince_rounds_mul_input_s2[27]), .B(
        prince_rounds_mul_s2_n68), .ZN(prince_rounds_mul_result_s2[19]) );
  XNOR2_X1 prince_rounds_mul_s2_U20 ( .A(prince_rounds_mul_input_s2[23]), .B(
        prince_rounds_mul_input_s2[19]), .ZN(prince_rounds_mul_s2_n68) );
  XNOR2_X1 prince_rounds_mul_s2_U19 ( .A(prince_rounds_mul_input_s2[22]), .B(
        prince_rounds_mul_s2_n67), .ZN(prince_rounds_mul_result_s2[18]) );
  XNOR2_X1 prince_rounds_mul_s2_U18 ( .A(prince_rounds_mul_input_s2[18]), .B(
        prince_rounds_mul_input_s2[30]), .ZN(prince_rounds_mul_s2_n67) );
  XNOR2_X1 prince_rounds_mul_s2_U17 ( .A(prince_rounds_mul_input_s2[29]), .B(
        prince_rounds_mul_s2_n70), .ZN(prince_rounds_mul_result_s2[17]) );
  XNOR2_X1 prince_rounds_mul_s2_U16 ( .A(prince_rounds_mul_input_s2[17]), .B(
        prince_rounds_mul_input_s2[25]), .ZN(prince_rounds_mul_s2_n70) );
  XNOR2_X1 prince_rounds_mul_s2_U15 ( .A(prince_rounds_mul_input_s2[20]), .B(
        prince_rounds_mul_s2_n71), .ZN(prince_rounds_mul_result_s2[16]) );
  XNOR2_X1 prince_rounds_mul_s2_U14 ( .A(prince_rounds_mul_input_s2[24]), .B(
        prince_rounds_mul_input_s2[28]), .ZN(prince_rounds_mul_s2_n71) );
  XNOR2_X1 prince_rounds_mul_s2_U13 ( .A(prince_rounds_mul_input_s2[3]), .B(
        prince_rounds_mul_s2_n65), .ZN(prince_rounds_mul_result_s2[15]) );
  XNOR2_X1 prince_rounds_mul_s2_U12 ( .A(prince_rounds_mul_input_s2[2]), .B(
        prince_rounds_mul_s2_n93), .ZN(prince_rounds_mul_result_s2[14]) );
  XNOR2_X1 prince_rounds_mul_s2_U11 ( .A(prince_rounds_mul_input_s2[6]), .B(
        prince_rounds_mul_input_s2[14]), .ZN(prince_rounds_mul_s2_n93) );
  XNOR2_X1 prince_rounds_mul_s2_U10 ( .A(prince_rounds_mul_input_s2[1]), .B(
        prince_rounds_mul_s2_n66), .ZN(prince_rounds_mul_result_s2[13]) );
  XNOR2_X1 prince_rounds_mul_s2_U9 ( .A(prince_rounds_mul_input_s2[13]), .B(
        prince_rounds_mul_input_s2[9]), .ZN(prince_rounds_mul_s2_n66) );
  XNOR2_X1 prince_rounds_mul_s2_U8 ( .A(prince_rounds_mul_input_s2[4]), .B(
        prince_rounds_mul_s2_n95), .ZN(prince_rounds_mul_result_s2[12]) );
  XNOR2_X1 prince_rounds_mul_s2_U7 ( .A(prince_rounds_mul_input_s2[8]), .B(
        prince_rounds_mul_input_s2[12]), .ZN(prince_rounds_mul_s2_n95) );
  XNOR2_X1 prince_rounds_mul_s2_U6 ( .A(prince_rounds_mul_input_s2[15]), .B(
        prince_rounds_mul_s2_n65), .ZN(prince_rounds_mul_result_s2[11]) );
  XNOR2_X1 prince_rounds_mul_s2_U5 ( .A(prince_rounds_mul_input_s2[11]), .B(
        prince_rounds_mul_input_s2[7]), .ZN(prince_rounds_mul_s2_n65) );
  XNOR2_X1 prince_rounds_mul_s2_U4 ( .A(prince_rounds_mul_input_s2[6]), .B(
        prince_rounds_mul_s2_n73), .ZN(prince_rounds_mul_result_s2[10]) );
  XNOR2_X1 prince_rounds_mul_s2_U3 ( .A(prince_rounds_mul_input_s2[10]), .B(
        prince_rounds_mul_input_s2[2]), .ZN(prince_rounds_mul_s2_n73) );
  XNOR2_X1 prince_rounds_mul_s2_U2 ( .A(prince_rounds_mul_input_s2[8]), .B(
        prince_rounds_mul_s2_n84), .ZN(prince_rounds_mul_result_s2[0]) );
  XNOR2_X1 prince_rounds_mul_s2_U1 ( .A(prince_rounds_mul_input_s2[0]), .B(
        prince_rounds_mul_input_s2[4]), .ZN(prince_rounds_mul_s2_n84) );
  XNOR2_X1 prince_rounds_mul_s3_U96 ( .A(prince_rounds_mul_input_s3[13]), .B(
        prince_rounds_mul_s3_n96), .ZN(prince_rounds_mul_result_s3[9]) );
  XNOR2_X1 prince_rounds_mul_s3_U95 ( .A(prince_rounds_mul_input_s3[0]), .B(
        prince_rounds_mul_s3_n95), .ZN(prince_rounds_mul_result_s3[8]) );
  XNOR2_X1 prince_rounds_mul_s3_U94 ( .A(prince_rounds_mul_input_s3[11]), .B(
        prince_rounds_mul_s3_n94), .ZN(prince_rounds_mul_result_s3[7]) );
  XNOR2_X1 prince_rounds_mul_s3_U93 ( .A(prince_rounds_mul_input_s3[10]), .B(
        prince_rounds_mul_s3_n93), .ZN(prince_rounds_mul_result_s3[6]) );
  XNOR2_X1 prince_rounds_mul_s3_U92 ( .A(prince_rounds_mul_input_s3[51]), .B(
        prince_rounds_mul_s3_n92), .ZN(prince_rounds_mul_result_s3[63]) );
  XNOR2_X1 prince_rounds_mul_s3_U91 ( .A(prince_rounds_mul_input_s3[50]), .B(
        prince_rounds_mul_s3_n91), .ZN(prince_rounds_mul_result_s3[62]) );
  XNOR2_X1 prince_rounds_mul_s3_U90 ( .A(prince_rounds_mul_input_s3[49]), .B(
        prince_rounds_mul_s3_n90), .ZN(prince_rounds_mul_result_s3[61]) );
  XNOR2_X1 prince_rounds_mul_s3_U89 ( .A(prince_rounds_mul_input_s3[52]), .B(
        prince_rounds_mul_s3_n89), .ZN(prince_rounds_mul_result_s3[60]) );
  XNOR2_X1 prince_rounds_mul_s3_U88 ( .A(prince_rounds_mul_input_s3[9]), .B(
        prince_rounds_mul_s3_n96), .ZN(prince_rounds_mul_result_s3[5]) );
  XNOR2_X1 prince_rounds_mul_s3_U87 ( .A(prince_rounds_mul_input_s3[1]), .B(
        prince_rounds_mul_input_s3[5]), .ZN(prince_rounds_mul_s3_n96) );
  XNOR2_X1 prince_rounds_mul_s3_U86 ( .A(prince_rounds_mul_input_s3[63]), .B(
        prince_rounds_mul_s3_n92), .ZN(prince_rounds_mul_result_s3[59]) );
  XNOR2_X1 prince_rounds_mul_s3_U85 ( .A(prince_rounds_mul_input_s3[55]), .B(
        prince_rounds_mul_input_s3[59]), .ZN(prince_rounds_mul_s3_n92) );
  XNOR2_X1 prince_rounds_mul_s3_U84 ( .A(prince_rounds_mul_input_s3[54]), .B(
        prince_rounds_mul_s3_n88), .ZN(prince_rounds_mul_result_s3[58]) );
  XNOR2_X1 prince_rounds_mul_s3_U83 ( .A(prince_rounds_mul_input_s3[61]), .B(
        prince_rounds_mul_s3_n87), .ZN(prince_rounds_mul_result_s3[57]) );
  XNOR2_X1 prince_rounds_mul_s3_U82 ( .A(prince_rounds_mul_input_s3[48]), .B(
        prince_rounds_mul_s3_n89), .ZN(prince_rounds_mul_result_s3[56]) );
  XNOR2_X1 prince_rounds_mul_s3_U81 ( .A(prince_rounds_mul_input_s3[56]), .B(
        prince_rounds_mul_input_s3[60]), .ZN(prince_rounds_mul_s3_n89) );
  XNOR2_X1 prince_rounds_mul_s3_U80 ( .A(prince_rounds_mul_input_s3[59]), .B(
        prince_rounds_mul_s3_n86), .ZN(prince_rounds_mul_result_s3[55]) );
  XNOR2_X1 prince_rounds_mul_s3_U79 ( .A(prince_rounds_mul_input_s3[58]), .B(
        prince_rounds_mul_s3_n91), .ZN(prince_rounds_mul_result_s3[54]) );
  XNOR2_X1 prince_rounds_mul_s3_U78 ( .A(prince_rounds_mul_input_s3[62]), .B(
        prince_rounds_mul_input_s3[54]), .ZN(prince_rounds_mul_s3_n91) );
  XNOR2_X1 prince_rounds_mul_s3_U77 ( .A(prince_rounds_mul_input_s3[57]), .B(
        prince_rounds_mul_s3_n87), .ZN(prince_rounds_mul_result_s3[53]) );
  XNOR2_X1 prince_rounds_mul_s3_U76 ( .A(prince_rounds_mul_input_s3[53]), .B(
        prince_rounds_mul_input_s3[49]), .ZN(prince_rounds_mul_s3_n87) );
  XNOR2_X1 prince_rounds_mul_s3_U75 ( .A(prince_rounds_mul_input_s3[60]), .B(
        prince_rounds_mul_s3_n85), .ZN(prince_rounds_mul_result_s3[52]) );
  XNOR2_X1 prince_rounds_mul_s3_U74 ( .A(prince_rounds_mul_input_s3[55]), .B(
        prince_rounds_mul_s3_n86), .ZN(prince_rounds_mul_result_s3[51]) );
  XNOR2_X1 prince_rounds_mul_s3_U73 ( .A(prince_rounds_mul_input_s3[51]), .B(
        prince_rounds_mul_input_s3[63]), .ZN(prince_rounds_mul_s3_n86) );
  XNOR2_X1 prince_rounds_mul_s3_U72 ( .A(prince_rounds_mul_input_s3[62]), .B(
        prince_rounds_mul_s3_n88), .ZN(prince_rounds_mul_result_s3[50]) );
  XNOR2_X1 prince_rounds_mul_s3_U71 ( .A(prince_rounds_mul_input_s3[50]), .B(
        prince_rounds_mul_input_s3[58]), .ZN(prince_rounds_mul_s3_n88) );
  XNOR2_X1 prince_rounds_mul_s3_U70 ( .A(prince_rounds_mul_input_s3[12]), .B(
        prince_rounds_mul_s3_n84), .ZN(prince_rounds_mul_result_s3[4]) );
  XNOR2_X1 prince_rounds_mul_s3_U69 ( .A(prince_rounds_mul_input_s3[53]), .B(
        prince_rounds_mul_s3_n90), .ZN(prince_rounds_mul_result_s3[49]) );
  XNOR2_X1 prince_rounds_mul_s3_U68 ( .A(prince_rounds_mul_input_s3[57]), .B(
        prince_rounds_mul_input_s3[61]), .ZN(prince_rounds_mul_s3_n90) );
  XNOR2_X1 prince_rounds_mul_s3_U67 ( .A(prince_rounds_mul_input_s3[56]), .B(
        prince_rounds_mul_s3_n85), .ZN(prince_rounds_mul_result_s3[48]) );
  XNOR2_X1 prince_rounds_mul_s3_U66 ( .A(prince_rounds_mul_input_s3[52]), .B(
        prince_rounds_mul_input_s3[48]), .ZN(prince_rounds_mul_s3_n85) );
  XNOR2_X1 prince_rounds_mul_s3_U65 ( .A(prince_rounds_mul_input_s3[39]), .B(
        prince_rounds_mul_s3_n83), .ZN(prince_rounds_mul_result_s3[47]) );
  XNOR2_X1 prince_rounds_mul_s3_U64 ( .A(prince_rounds_mul_input_s3[34]), .B(
        prince_rounds_mul_s3_n82), .ZN(prince_rounds_mul_result_s3[46]) );
  XNOR2_X1 prince_rounds_mul_s3_U63 ( .A(prince_rounds_mul_input_s3[33]), .B(
        prince_rounds_mul_s3_n81), .ZN(prince_rounds_mul_result_s3[45]) );
  XNOR2_X1 prince_rounds_mul_s3_U62 ( .A(prince_rounds_mul_input_s3[32]), .B(
        prince_rounds_mul_s3_n80), .ZN(prince_rounds_mul_result_s3[44]) );
  XNOR2_X1 prince_rounds_mul_s3_U61 ( .A(prince_rounds_mul_input_s3[35]), .B(
        prince_rounds_mul_s3_n83), .ZN(prince_rounds_mul_result_s3[43]) );
  XNOR2_X1 prince_rounds_mul_s3_U60 ( .A(prince_rounds_mul_input_s3[43]), .B(
        prince_rounds_mul_input_s3[47]), .ZN(prince_rounds_mul_s3_n83) );
  XNOR2_X1 prince_rounds_mul_s3_U59 ( .A(prince_rounds_mul_input_s3[46]), .B(
        prince_rounds_mul_s3_n82), .ZN(prince_rounds_mul_result_s3[42]) );
  XNOR2_X1 prince_rounds_mul_s3_U58 ( .A(prince_rounds_mul_input_s3[38]), .B(
        prince_rounds_mul_input_s3[42]), .ZN(prince_rounds_mul_s3_n82) );
  XNOR2_X1 prince_rounds_mul_s3_U57 ( .A(prince_rounds_mul_input_s3[37]), .B(
        prince_rounds_mul_s3_n79), .ZN(prince_rounds_mul_result_s3[41]) );
  XNOR2_X1 prince_rounds_mul_s3_U56 ( .A(prince_rounds_mul_input_s3[44]), .B(
        prince_rounds_mul_s3_n78), .ZN(prince_rounds_mul_result_s3[40]) );
  XNOR2_X1 prince_rounds_mul_s3_U55 ( .A(prince_rounds_mul_input_s3[7]), .B(
        prince_rounds_mul_s3_n94), .ZN(prince_rounds_mul_result_s3[3]) );
  XNOR2_X1 prince_rounds_mul_s3_U54 ( .A(prince_rounds_mul_input_s3[15]), .B(
        prince_rounds_mul_input_s3[3]), .ZN(prince_rounds_mul_s3_n94) );
  XNOR2_X1 prince_rounds_mul_s3_U53 ( .A(prince_rounds_mul_input_s3[47]), .B(
        prince_rounds_mul_s3_n77), .ZN(prince_rounds_mul_result_s3[39]) );
  XNOR2_X1 prince_rounds_mul_s3_U52 ( .A(prince_rounds_mul_input_s3[42]), .B(
        prince_rounds_mul_s3_n76), .ZN(prince_rounds_mul_result_s3[38]) );
  XNOR2_X1 prince_rounds_mul_s3_U51 ( .A(prince_rounds_mul_input_s3[41]), .B(
        prince_rounds_mul_s3_n81), .ZN(prince_rounds_mul_result_s3[37]) );
  XNOR2_X1 prince_rounds_mul_s3_U50 ( .A(prince_rounds_mul_input_s3[45]), .B(
        prince_rounds_mul_input_s3[37]), .ZN(prince_rounds_mul_s3_n81) );
  XNOR2_X1 prince_rounds_mul_s3_U49 ( .A(prince_rounds_mul_input_s3[40]), .B(
        prince_rounds_mul_s3_n78), .ZN(prince_rounds_mul_result_s3[36]) );
  XNOR2_X1 prince_rounds_mul_s3_U48 ( .A(prince_rounds_mul_input_s3[36]), .B(
        prince_rounds_mul_input_s3[32]), .ZN(prince_rounds_mul_s3_n78) );
  XNOR2_X1 prince_rounds_mul_s3_U47 ( .A(prince_rounds_mul_input_s3[43]), .B(
        prince_rounds_mul_s3_n77), .ZN(prince_rounds_mul_result_s3[35]) );
  XNOR2_X1 prince_rounds_mul_s3_U46 ( .A(prince_rounds_mul_input_s3[39]), .B(
        prince_rounds_mul_input_s3[35]), .ZN(prince_rounds_mul_s3_n77) );
  XNOR2_X1 prince_rounds_mul_s3_U45 ( .A(prince_rounds_mul_input_s3[38]), .B(
        prince_rounds_mul_s3_n76), .ZN(prince_rounds_mul_result_s3[34]) );
  XNOR2_X1 prince_rounds_mul_s3_U44 ( .A(prince_rounds_mul_input_s3[34]), .B(
        prince_rounds_mul_input_s3[46]), .ZN(prince_rounds_mul_s3_n76) );
  XNOR2_X1 prince_rounds_mul_s3_U43 ( .A(prince_rounds_mul_input_s3[45]), .B(
        prince_rounds_mul_s3_n79), .ZN(prince_rounds_mul_result_s3[33]) );
  XNOR2_X1 prince_rounds_mul_s3_U42 ( .A(prince_rounds_mul_input_s3[33]), .B(
        prince_rounds_mul_input_s3[41]), .ZN(prince_rounds_mul_s3_n79) );
  XNOR2_X1 prince_rounds_mul_s3_U41 ( .A(prince_rounds_mul_input_s3[36]), .B(
        prince_rounds_mul_s3_n80), .ZN(prince_rounds_mul_result_s3[32]) );
  XNOR2_X1 prince_rounds_mul_s3_U40 ( .A(prince_rounds_mul_input_s3[40]), .B(
        prince_rounds_mul_input_s3[44]), .ZN(prince_rounds_mul_s3_n80) );
  XNOR2_X1 prince_rounds_mul_s3_U39 ( .A(prince_rounds_mul_input_s3[23]), .B(
        prince_rounds_mul_s3_n75), .ZN(prince_rounds_mul_result_s3[31]) );
  XNOR2_X1 prince_rounds_mul_s3_U38 ( .A(prince_rounds_mul_input_s3[18]), .B(
        prince_rounds_mul_s3_n74), .ZN(prince_rounds_mul_result_s3[30]) );
  XNOR2_X1 prince_rounds_mul_s3_U37 ( .A(prince_rounds_mul_input_s3[14]), .B(
        prince_rounds_mul_s3_n73), .ZN(prince_rounds_mul_result_s3[2]) );
  XNOR2_X1 prince_rounds_mul_s3_U36 ( .A(prince_rounds_mul_input_s3[17]), .B(
        prince_rounds_mul_s3_n72), .ZN(prince_rounds_mul_result_s3[29]) );
  XNOR2_X1 prince_rounds_mul_s3_U35 ( .A(prince_rounds_mul_input_s3[16]), .B(
        prince_rounds_mul_s3_n71), .ZN(prince_rounds_mul_result_s3[28]) );
  XNOR2_X1 prince_rounds_mul_s3_U34 ( .A(prince_rounds_mul_input_s3[19]), .B(
        prince_rounds_mul_s3_n75), .ZN(prince_rounds_mul_result_s3[27]) );
  XNOR2_X1 prince_rounds_mul_s3_U33 ( .A(prince_rounds_mul_input_s3[27]), .B(
        prince_rounds_mul_input_s3[31]), .ZN(prince_rounds_mul_s3_n75) );
  XNOR2_X1 prince_rounds_mul_s3_U32 ( .A(prince_rounds_mul_input_s3[30]), .B(
        prince_rounds_mul_s3_n74), .ZN(prince_rounds_mul_result_s3[26]) );
  XNOR2_X1 prince_rounds_mul_s3_U31 ( .A(prince_rounds_mul_input_s3[22]), .B(
        prince_rounds_mul_input_s3[26]), .ZN(prince_rounds_mul_s3_n74) );
  XNOR2_X1 prince_rounds_mul_s3_U30 ( .A(prince_rounds_mul_input_s3[21]), .B(
        prince_rounds_mul_s3_n70), .ZN(prince_rounds_mul_result_s3[25]) );
  XNOR2_X1 prince_rounds_mul_s3_U29 ( .A(prince_rounds_mul_input_s3[28]), .B(
        prince_rounds_mul_s3_n69), .ZN(prince_rounds_mul_result_s3[24]) );
  XNOR2_X1 prince_rounds_mul_s3_U28 ( .A(prince_rounds_mul_input_s3[31]), .B(
        prince_rounds_mul_s3_n68), .ZN(prince_rounds_mul_result_s3[23]) );
  XNOR2_X1 prince_rounds_mul_s3_U27 ( .A(prince_rounds_mul_input_s3[26]), .B(
        prince_rounds_mul_s3_n67), .ZN(prince_rounds_mul_result_s3[22]) );
  XNOR2_X1 prince_rounds_mul_s3_U26 ( .A(prince_rounds_mul_input_s3[25]), .B(
        prince_rounds_mul_s3_n72), .ZN(prince_rounds_mul_result_s3[21]) );
  XNOR2_X1 prince_rounds_mul_s3_U25 ( .A(prince_rounds_mul_input_s3[29]), .B(
        prince_rounds_mul_input_s3[21]), .ZN(prince_rounds_mul_s3_n72) );
  XNOR2_X1 prince_rounds_mul_s3_U24 ( .A(prince_rounds_mul_input_s3[24]), .B(
        prince_rounds_mul_s3_n69), .ZN(prince_rounds_mul_result_s3[20]) );
  XNOR2_X1 prince_rounds_mul_s3_U23 ( .A(prince_rounds_mul_input_s3[20]), .B(
        prince_rounds_mul_input_s3[16]), .ZN(prince_rounds_mul_s3_n69) );
  XNOR2_X1 prince_rounds_mul_s3_U22 ( .A(prince_rounds_mul_input_s3[5]), .B(
        prince_rounds_mul_s3_n66), .ZN(prince_rounds_mul_result_s3[1]) );
  XNOR2_X1 prince_rounds_mul_s3_U21 ( .A(prince_rounds_mul_input_s3[27]), .B(
        prince_rounds_mul_s3_n68), .ZN(prince_rounds_mul_result_s3[19]) );
  XNOR2_X1 prince_rounds_mul_s3_U20 ( .A(prince_rounds_mul_input_s3[23]), .B(
        prince_rounds_mul_input_s3[19]), .ZN(prince_rounds_mul_s3_n68) );
  XNOR2_X1 prince_rounds_mul_s3_U19 ( .A(prince_rounds_mul_input_s3[22]), .B(
        prince_rounds_mul_s3_n67), .ZN(prince_rounds_mul_result_s3[18]) );
  XNOR2_X1 prince_rounds_mul_s3_U18 ( .A(prince_rounds_mul_input_s3[18]), .B(
        prince_rounds_mul_input_s3[30]), .ZN(prince_rounds_mul_s3_n67) );
  XNOR2_X1 prince_rounds_mul_s3_U17 ( .A(prince_rounds_mul_input_s3[29]), .B(
        prince_rounds_mul_s3_n70), .ZN(prince_rounds_mul_result_s3[17]) );
  XNOR2_X1 prince_rounds_mul_s3_U16 ( .A(prince_rounds_mul_input_s3[17]), .B(
        prince_rounds_mul_input_s3[25]), .ZN(prince_rounds_mul_s3_n70) );
  XNOR2_X1 prince_rounds_mul_s3_U15 ( .A(prince_rounds_mul_input_s3[20]), .B(
        prince_rounds_mul_s3_n71), .ZN(prince_rounds_mul_result_s3[16]) );
  XNOR2_X1 prince_rounds_mul_s3_U14 ( .A(prince_rounds_mul_input_s3[24]), .B(
        prince_rounds_mul_input_s3[28]), .ZN(prince_rounds_mul_s3_n71) );
  XNOR2_X1 prince_rounds_mul_s3_U13 ( .A(prince_rounds_mul_input_s3[3]), .B(
        prince_rounds_mul_s3_n65), .ZN(prince_rounds_mul_result_s3[15]) );
  XNOR2_X1 prince_rounds_mul_s3_U12 ( .A(prince_rounds_mul_input_s3[2]), .B(
        prince_rounds_mul_s3_n93), .ZN(prince_rounds_mul_result_s3[14]) );
  XNOR2_X1 prince_rounds_mul_s3_U11 ( .A(prince_rounds_mul_input_s3[6]), .B(
        prince_rounds_mul_input_s3[14]), .ZN(prince_rounds_mul_s3_n93) );
  XNOR2_X1 prince_rounds_mul_s3_U10 ( .A(prince_rounds_mul_input_s3[1]), .B(
        prince_rounds_mul_s3_n66), .ZN(prince_rounds_mul_result_s3[13]) );
  XNOR2_X1 prince_rounds_mul_s3_U9 ( .A(prince_rounds_mul_input_s3[13]), .B(
        prince_rounds_mul_input_s3[9]), .ZN(prince_rounds_mul_s3_n66) );
  XNOR2_X1 prince_rounds_mul_s3_U8 ( .A(prince_rounds_mul_input_s3[4]), .B(
        prince_rounds_mul_s3_n95), .ZN(prince_rounds_mul_result_s3[12]) );
  XNOR2_X1 prince_rounds_mul_s3_U7 ( .A(prince_rounds_mul_input_s3[8]), .B(
        prince_rounds_mul_input_s3[12]), .ZN(prince_rounds_mul_s3_n95) );
  XNOR2_X1 prince_rounds_mul_s3_U6 ( .A(prince_rounds_mul_input_s3[15]), .B(
        prince_rounds_mul_s3_n65), .ZN(prince_rounds_mul_result_s3[11]) );
  XNOR2_X1 prince_rounds_mul_s3_U5 ( .A(prince_rounds_mul_input_s3[11]), .B(
        prince_rounds_mul_input_s3[7]), .ZN(prince_rounds_mul_s3_n65) );
  XNOR2_X1 prince_rounds_mul_s3_U4 ( .A(prince_rounds_mul_input_s3[6]), .B(
        prince_rounds_mul_s3_n73), .ZN(prince_rounds_mul_result_s3[10]) );
  XNOR2_X1 prince_rounds_mul_s3_U3 ( .A(prince_rounds_mul_input_s3[10]), .B(
        prince_rounds_mul_input_s3[2]), .ZN(prince_rounds_mul_s3_n73) );
  XNOR2_X1 prince_rounds_mul_s3_U2 ( .A(prince_rounds_mul_input_s3[8]), .B(
        prince_rounds_mul_s3_n84), .ZN(prince_rounds_mul_result_s3[0]) );
  XNOR2_X1 prince_rounds_mul_s3_U1 ( .A(prince_rounds_mul_input_s3[0]), .B(
        prince_rounds_mul_input_s3[4]), .ZN(prince_rounds_mul_s3_n84) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_0_0_U2 ( .A(
        prince_AddKeyOut1_XORInst_0_0_n3), .B(prince_selected_Key1_0_), .ZN(
        output_s1[0]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_0_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[0]), .ZN(prince_AddKeyOut1_XORInst_0_0_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_0_1_U2 ( .A(
        prince_AddKeyOut1_XORInst_0_1_n3), .B(prince_selected_Key1_1_), .ZN(
        output_s1[1]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_0_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[1]), .ZN(prince_AddKeyOut1_XORInst_0_1_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_0_2_U2 ( .A(
        prince_AddKeyOut1_XORInst_0_2_n3), .B(prince_selected_Key1_2_), .ZN(
        output_s1[2]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_0_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[2]), .ZN(prince_AddKeyOut1_XORInst_0_2_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_0_3_U2 ( .A(
        prince_AddKeyOut1_XORInst_0_3_n3), .B(prince_selected_Key1_3_), .ZN(
        output_s1[3]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_0_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[3]), .ZN(prince_AddKeyOut1_XORInst_0_3_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_1_0_U2 ( .A(
        prince_AddKeyOut1_XORInst_1_0_n3), .B(prince_selected_Key1_4_), .ZN(
        output_s1[4]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_1_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[4]), .ZN(prince_AddKeyOut1_XORInst_1_0_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_1_1_U2 ( .A(
        prince_AddKeyOut1_XORInst_1_1_n3), .B(prince_selected_Key1_5_), .ZN(
        output_s1[5]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_1_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[5]), .ZN(prince_AddKeyOut1_XORInst_1_1_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_1_2_U2 ( .A(
        prince_AddKeyOut1_XORInst_1_2_n3), .B(prince_selected_Key1_6_), .ZN(
        output_s1[6]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_1_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[6]), .ZN(prince_AddKeyOut1_XORInst_1_2_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_1_3_U2 ( .A(
        prince_AddKeyOut1_XORInst_1_3_n3), .B(prince_selected_Key1_7_), .ZN(
        output_s1[7]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_1_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[7]), .ZN(prince_AddKeyOut1_XORInst_1_3_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_2_0_U2 ( .A(
        prince_AddKeyOut1_XORInst_2_0_n3), .B(prince_selected_Key1_8_), .ZN(
        output_s1[8]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_2_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[8]), .ZN(prince_AddKeyOut1_XORInst_2_0_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_2_1_U2 ( .A(
        prince_AddKeyOut1_XORInst_2_1_n3), .B(prince_selected_Key1_9_), .ZN(
        output_s1[9]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_2_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[9]), .ZN(prince_AddKeyOut1_XORInst_2_1_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_2_2_U2 ( .A(
        prince_AddKeyOut1_XORInst_2_2_n3), .B(prince_selected_Key1_10_), .ZN(
        output_s1[10]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_2_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[10]), .ZN(prince_AddKeyOut1_XORInst_2_2_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_2_3_U2 ( .A(
        prince_AddKeyOut1_XORInst_2_3_n3), .B(prince_selected_Key1_11_), .ZN(
        output_s1[11]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_2_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[11]), .ZN(prince_AddKeyOut1_XORInst_2_3_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_3_0_U2 ( .A(
        prince_AddKeyOut1_XORInst_3_0_n3), .B(prince_selected_Key1_12_), .ZN(
        output_s1[12]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_3_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[12]), .ZN(prince_AddKeyOut1_XORInst_3_0_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_3_1_U2 ( .A(
        prince_AddKeyOut1_XORInst_3_1_n3), .B(prince_selected_Key1_13_), .ZN(
        output_s1[13]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_3_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[13]), .ZN(prince_AddKeyOut1_XORInst_3_1_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_3_2_U2 ( .A(
        prince_AddKeyOut1_XORInst_3_2_n3), .B(prince_selected_Key1_14_), .ZN(
        output_s1[14]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_3_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[14]), .ZN(prince_AddKeyOut1_XORInst_3_2_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_3_3_U2 ( .A(
        prince_AddKeyOut1_XORInst_3_3_n3), .B(prince_selected_Key1_15_), .ZN(
        output_s1[15]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_3_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[15]), .ZN(prince_AddKeyOut1_XORInst_3_3_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_4_0_U2 ( .A(
        prince_AddKeyOut1_XORInst_4_0_n3), .B(prince_selected_Key1_16_), .ZN(
        output_s1[16]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_4_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[16]), .ZN(prince_AddKeyOut1_XORInst_4_0_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_4_1_U2 ( .A(
        prince_AddKeyOut1_XORInst_4_1_n3), .B(prince_selected_Key1_17_), .ZN(
        output_s1[17]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_4_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[17]), .ZN(prince_AddKeyOut1_XORInst_4_1_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_4_2_U2 ( .A(
        prince_AddKeyOut1_XORInst_4_2_n3), .B(prince_selected_Key1_18_), .ZN(
        output_s1[18]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_4_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[18]), .ZN(prince_AddKeyOut1_XORInst_4_2_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_4_3_U2 ( .A(
        prince_AddKeyOut1_XORInst_4_3_n3), .B(prince_selected_Key1_19_), .ZN(
        output_s1[19]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_4_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[19]), .ZN(prince_AddKeyOut1_XORInst_4_3_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_5_0_U2 ( .A(
        prince_AddKeyOut1_XORInst_5_0_n3), .B(prince_selected_Key1_20_), .ZN(
        output_s1[20]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_5_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[20]), .ZN(prince_AddKeyOut1_XORInst_5_0_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_5_1_U2 ( .A(
        prince_AddKeyOut1_XORInst_5_1_n3), .B(prince_selected_Key1_21_), .ZN(
        output_s1[21]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_5_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[21]), .ZN(prince_AddKeyOut1_XORInst_5_1_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_5_2_U2 ( .A(
        prince_AddKeyOut1_XORInst_5_2_n3), .B(prince_selected_Key1_22_), .ZN(
        output_s1[22]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_5_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[22]), .ZN(prince_AddKeyOut1_XORInst_5_2_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_5_3_U2 ( .A(
        prince_AddKeyOut1_XORInst_5_3_n3), .B(prince_selected_Key1_23_), .ZN(
        output_s1[23]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_5_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[23]), .ZN(prince_AddKeyOut1_XORInst_5_3_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_6_0_U2 ( .A(
        prince_AddKeyOut1_XORInst_6_0_n3), .B(prince_selected_Key1_24_), .ZN(
        output_s1[24]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_6_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[24]), .ZN(prince_AddKeyOut1_XORInst_6_0_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_6_1_U2 ( .A(
        prince_AddKeyOut1_XORInst_6_1_n3), .B(prince_selected_Key1_25_), .ZN(
        output_s1[25]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_6_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[25]), .ZN(prince_AddKeyOut1_XORInst_6_1_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_6_2_U2 ( .A(
        prince_AddKeyOut1_XORInst_6_2_n3), .B(prince_selected_Key1_26_), .ZN(
        output_s1[26]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_6_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[26]), .ZN(prince_AddKeyOut1_XORInst_6_2_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_6_3_U2 ( .A(
        prince_AddKeyOut1_XORInst_6_3_n3), .B(prince_selected_Key1_27_), .ZN(
        output_s1[27]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_6_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[27]), .ZN(prince_AddKeyOut1_XORInst_6_3_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_7_0_U2 ( .A(
        prince_AddKeyOut1_XORInst_7_0_n3), .B(prince_selected_Key1_28_), .ZN(
        output_s1[28]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_7_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[28]), .ZN(prince_AddKeyOut1_XORInst_7_0_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_7_1_U2 ( .A(
        prince_AddKeyOut1_XORInst_7_1_n3), .B(prince_selected_Key1_29_), .ZN(
        output_s1[29]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_7_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[29]), .ZN(prince_AddKeyOut1_XORInst_7_1_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_7_2_U2 ( .A(
        prince_AddKeyOut1_XORInst_7_2_n3), .B(prince_selected_Key1_30_), .ZN(
        output_s1[30]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_7_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[30]), .ZN(prince_AddKeyOut1_XORInst_7_2_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_7_3_U2 ( .A(
        prince_AddKeyOut1_XORInst_7_3_n3), .B(prince_selected_Key1_31_), .ZN(
        output_s1[31]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_7_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[31]), .ZN(prince_AddKeyOut1_XORInst_7_3_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_8_0_U2 ( .A(
        prince_AddKeyOut1_XORInst_8_0_n3), .B(prince_selected_Key1_32_), .ZN(
        output_s1[32]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_8_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[32]), .ZN(prince_AddKeyOut1_XORInst_8_0_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_8_1_U2 ( .A(
        prince_AddKeyOut1_XORInst_8_1_n3), .B(prince_selected_Key1_33_), .ZN(
        output_s1[33]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_8_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[33]), .ZN(prince_AddKeyOut1_XORInst_8_1_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_8_2_U2 ( .A(
        prince_AddKeyOut1_XORInst_8_2_n3), .B(prince_selected_Key1_34_), .ZN(
        output_s1[34]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_8_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[34]), .ZN(prince_AddKeyOut1_XORInst_8_2_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_8_3_U2 ( .A(
        prince_AddKeyOut1_XORInst_8_3_n3), .B(prince_selected_Key1_35_), .ZN(
        output_s1[35]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_8_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[35]), .ZN(prince_AddKeyOut1_XORInst_8_3_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_9_0_U2 ( .A(
        prince_AddKeyOut1_XORInst_9_0_n3), .B(prince_selected_Key1_36_), .ZN(
        output_s1[36]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_9_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[36]), .ZN(prince_AddKeyOut1_XORInst_9_0_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_9_1_U2 ( .A(
        prince_AddKeyOut1_XORInst_9_1_n3), .B(prince_selected_Key1_37_), .ZN(
        output_s1[37]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_9_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[37]), .ZN(prince_AddKeyOut1_XORInst_9_1_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_9_2_U2 ( .A(
        prince_AddKeyOut1_XORInst_9_2_n3), .B(prince_selected_Key1_38_), .ZN(
        output_s1[38]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_9_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[38]), .ZN(prince_AddKeyOut1_XORInst_9_2_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_9_3_U2 ( .A(
        prince_AddKeyOut1_XORInst_9_3_n3), .B(prince_selected_Key1_39_), .ZN(
        output_s1[39]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_9_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[39]), .ZN(prince_AddKeyOut1_XORInst_9_3_n3) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_10_0_U2 ( .A(
        prince_AddKeyOut1_XORInst_10_0_n3), .B(prince_selected_Key1_40_), .ZN(
        output_s1[40]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_10_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[40]), .ZN(prince_AddKeyOut1_XORInst_10_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_10_1_U2 ( .A(
        prince_AddKeyOut1_XORInst_10_1_n3), .B(prince_selected_Key1_41_), .ZN(
        output_s1[41]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_10_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[41]), .ZN(prince_AddKeyOut1_XORInst_10_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_10_2_U2 ( .A(
        prince_AddKeyOut1_XORInst_10_2_n3), .B(prince_selected_Key1_42_), .ZN(
        output_s1[42]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_10_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[42]), .ZN(prince_AddKeyOut1_XORInst_10_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_10_3_U2 ( .A(
        prince_AddKeyOut1_XORInst_10_3_n3), .B(prince_selected_Key1_43_), .ZN(
        output_s1[43]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_10_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[43]), .ZN(prince_AddKeyOut1_XORInst_10_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_11_0_U2 ( .A(
        prince_AddKeyOut1_XORInst_11_0_n3), .B(prince_selected_Key1_44_), .ZN(
        output_s1[44]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_11_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[44]), .ZN(prince_AddKeyOut1_XORInst_11_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_11_1_U2 ( .A(
        prince_AddKeyOut1_XORInst_11_1_n3), .B(prince_selected_Key1_45_), .ZN(
        output_s1[45]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_11_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[45]), .ZN(prince_AddKeyOut1_XORInst_11_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_11_2_U2 ( .A(
        prince_AddKeyOut1_XORInst_11_2_n3), .B(prince_selected_Key1_46_), .ZN(
        output_s1[46]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_11_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[46]), .ZN(prince_AddKeyOut1_XORInst_11_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_11_3_U2 ( .A(
        prince_AddKeyOut1_XORInst_11_3_n3), .B(prince_selected_Key1_47_), .ZN(
        output_s1[47]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_11_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[47]), .ZN(prince_AddKeyOut1_XORInst_11_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_12_0_U2 ( .A(
        prince_AddKeyOut1_XORInst_12_0_n3), .B(prince_selected_Key1_48_), .ZN(
        output_s1[48]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_12_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[48]), .ZN(prince_AddKeyOut1_XORInst_12_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_12_1_U2 ( .A(
        prince_AddKeyOut1_XORInst_12_1_n3), .B(prince_selected_Key1_49_), .ZN(
        output_s1[49]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_12_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[49]), .ZN(prince_AddKeyOut1_XORInst_12_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_12_2_U2 ( .A(
        prince_AddKeyOut1_XORInst_12_2_n3), .B(prince_selected_Key1_50_), .ZN(
        output_s1[50]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_12_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[50]), .ZN(prince_AddKeyOut1_XORInst_12_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_12_3_U2 ( .A(
        prince_AddKeyOut1_XORInst_12_3_n3), .B(prince_selected_Key1_51_), .ZN(
        output_s1[51]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_12_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[51]), .ZN(prince_AddKeyOut1_XORInst_12_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_13_0_U2 ( .A(
        prince_AddKeyOut1_XORInst_13_0_n3), .B(prince_selected_Key1_52_), .ZN(
        output_s1[52]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_13_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[52]), .ZN(prince_AddKeyOut1_XORInst_13_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_13_1_U2 ( .A(
        prince_AddKeyOut1_XORInst_13_1_n3), .B(prince_selected_Key1_53_), .ZN(
        output_s1[53]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_13_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[53]), .ZN(prince_AddKeyOut1_XORInst_13_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_13_2_U2 ( .A(
        prince_AddKeyOut1_XORInst_13_2_n3), .B(prince_selected_Key1_54_), .ZN(
        output_s1[54]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_13_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[54]), .ZN(prince_AddKeyOut1_XORInst_13_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_13_3_U2 ( .A(
        prince_AddKeyOut1_XORInst_13_3_n3), .B(prince_selected_Key1_55_), .ZN(
        output_s1[55]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_13_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[55]), .ZN(prince_AddKeyOut1_XORInst_13_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_14_0_U2 ( .A(
        prince_AddKeyOut1_XORInst_14_0_n3), .B(prince_selected_Key1_56_), .ZN(
        output_s1[56]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_14_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[56]), .ZN(prince_AddKeyOut1_XORInst_14_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_14_1_U2 ( .A(
        prince_AddKeyOut1_XORInst_14_1_n3), .B(prince_selected_Key1_57_), .ZN(
        output_s1[57]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_14_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[57]), .ZN(prince_AddKeyOut1_XORInst_14_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_14_2_U2 ( .A(
        prince_AddKeyOut1_XORInst_14_2_n3), .B(prince_selected_Key1_58_), .ZN(
        output_s1[58]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_14_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[58]), .ZN(prince_AddKeyOut1_XORInst_14_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_14_3_U2 ( .A(
        prince_AddKeyOut1_XORInst_14_3_n3), .B(prince_selected_Key1_59_), .ZN(
        output_s1[59]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_14_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[59]), .ZN(prince_AddKeyOut1_XORInst_14_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_15_0_U2 ( .A(
        prince_AddKeyOut1_XORInst_15_0_n3), .B(prince_selected_Key1_60_), .ZN(
        output_s1[60]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_15_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[60]), .ZN(prince_AddKeyOut1_XORInst_15_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_15_1_U2 ( .A(
        prince_AddKeyOut1_XORInst_15_1_n3), .B(prince_selected_Key1_61_), .ZN(
        output_s1[61]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_15_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[61]), .ZN(prince_AddKeyOut1_XORInst_15_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_15_2_U2 ( .A(
        prince_AddKeyOut1_XORInst_15_2_n3), .B(prince_selected_Key1_62_), .ZN(
        output_s1[62]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_15_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[62]), .ZN(prince_AddKeyOut1_XORInst_15_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut1_XORInst_15_3_U2 ( .A(
        prince_AddKeyOut1_XORInst_15_3_n3), .B(prince_selected_Key1_63_), .ZN(
        output_s1[63]) );
  XNOR2_X1 prince_AddKeyOut1_XORInst_15_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s1[63]), .ZN(prince_AddKeyOut1_XORInst_15_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_0_0_U2 ( .A(
        prince_AddKeyOut2_XORInst_0_0_n3), .B(prince_selected_Key2_0_), .ZN(
        output_s2[0]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_0_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[0]), .ZN(prince_AddKeyOut2_XORInst_0_0_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_0_1_U2 ( .A(
        prince_AddKeyOut2_XORInst_0_1_n3), .B(prince_selected_Key2_1_), .ZN(
        output_s2[1]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_0_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[1]), .ZN(prince_AddKeyOut2_XORInst_0_1_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_0_2_U2 ( .A(
        prince_AddKeyOut2_XORInst_0_2_n3), .B(prince_selected_Key2_2_), .ZN(
        output_s2[2]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_0_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[2]), .ZN(prince_AddKeyOut2_XORInst_0_2_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_0_3_U2 ( .A(
        prince_AddKeyOut2_XORInst_0_3_n3), .B(prince_selected_Key2_3_), .ZN(
        output_s2[3]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_0_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[3]), .ZN(prince_AddKeyOut2_XORInst_0_3_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_1_0_U2 ( .A(
        prince_AddKeyOut2_XORInst_1_0_n3), .B(prince_selected_Key2_4_), .ZN(
        output_s2[4]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_1_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[4]), .ZN(prince_AddKeyOut2_XORInst_1_0_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_1_1_U2 ( .A(
        prince_AddKeyOut2_XORInst_1_1_n3), .B(prince_selected_Key2_5_), .ZN(
        output_s2[5]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_1_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[5]), .ZN(prince_AddKeyOut2_XORInst_1_1_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_1_2_U2 ( .A(
        prince_AddKeyOut2_XORInst_1_2_n3), .B(prince_selected_Key2_6_), .ZN(
        output_s2[6]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_1_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[6]), .ZN(prince_AddKeyOut2_XORInst_1_2_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_1_3_U2 ( .A(
        prince_AddKeyOut2_XORInst_1_3_n3), .B(prince_selected_Key2_7_), .ZN(
        output_s2[7]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_1_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[7]), .ZN(prince_AddKeyOut2_XORInst_1_3_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_2_0_U2 ( .A(
        prince_AddKeyOut2_XORInst_2_0_n3), .B(prince_selected_Key2_8_), .ZN(
        output_s2[8]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_2_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[8]), .ZN(prince_AddKeyOut2_XORInst_2_0_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_2_1_U2 ( .A(
        prince_AddKeyOut2_XORInst_2_1_n3), .B(prince_selected_Key2_9_), .ZN(
        output_s2[9]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_2_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[9]), .ZN(prince_AddKeyOut2_XORInst_2_1_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_2_2_U2 ( .A(
        prince_AddKeyOut2_XORInst_2_2_n3), .B(prince_selected_Key2_10_), .ZN(
        output_s2[10]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_2_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[10]), .ZN(prince_AddKeyOut2_XORInst_2_2_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_2_3_U2 ( .A(
        prince_AddKeyOut2_XORInst_2_3_n3), .B(prince_selected_Key2_11_), .ZN(
        output_s2[11]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_2_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[11]), .ZN(prince_AddKeyOut2_XORInst_2_3_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_3_0_U2 ( .A(
        prince_AddKeyOut2_XORInst_3_0_n3), .B(prince_selected_Key2_12_), .ZN(
        output_s2[12]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_3_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[12]), .ZN(prince_AddKeyOut2_XORInst_3_0_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_3_1_U2 ( .A(
        prince_AddKeyOut2_XORInst_3_1_n3), .B(prince_selected_Key2_13_), .ZN(
        output_s2[13]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_3_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[13]), .ZN(prince_AddKeyOut2_XORInst_3_1_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_3_2_U2 ( .A(
        prince_AddKeyOut2_XORInst_3_2_n3), .B(prince_selected_Key2_14_), .ZN(
        output_s2[14]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_3_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[14]), .ZN(prince_AddKeyOut2_XORInst_3_2_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_3_3_U2 ( .A(
        prince_AddKeyOut2_XORInst_3_3_n3), .B(prince_selected_Key2_15_), .ZN(
        output_s2[15]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_3_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[15]), .ZN(prince_AddKeyOut2_XORInst_3_3_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_4_0_U2 ( .A(
        prince_AddKeyOut2_XORInst_4_0_n3), .B(prince_selected_Key2_16_), .ZN(
        output_s2[16]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_4_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[16]), .ZN(prince_AddKeyOut2_XORInst_4_0_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_4_1_U2 ( .A(
        prince_AddKeyOut2_XORInst_4_1_n3), .B(prince_selected_Key2_17_), .ZN(
        output_s2[17]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_4_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[17]), .ZN(prince_AddKeyOut2_XORInst_4_1_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_4_2_U2 ( .A(
        prince_AddKeyOut2_XORInst_4_2_n3), .B(prince_selected_Key2_18_), .ZN(
        output_s2[18]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_4_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[18]), .ZN(prince_AddKeyOut2_XORInst_4_2_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_4_3_U2 ( .A(
        prince_AddKeyOut2_XORInst_4_3_n3), .B(prince_selected_Key2_19_), .ZN(
        output_s2[19]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_4_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[19]), .ZN(prince_AddKeyOut2_XORInst_4_3_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_5_0_U2 ( .A(
        prince_AddKeyOut2_XORInst_5_0_n3), .B(prince_selected_Key2_20_), .ZN(
        output_s2[20]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_5_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[20]), .ZN(prince_AddKeyOut2_XORInst_5_0_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_5_1_U2 ( .A(
        prince_AddKeyOut2_XORInst_5_1_n3), .B(prince_selected_Key2_21_), .ZN(
        output_s2[21]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_5_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[21]), .ZN(prince_AddKeyOut2_XORInst_5_1_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_5_2_U2 ( .A(
        prince_AddKeyOut2_XORInst_5_2_n3), .B(prince_selected_Key2_22_), .ZN(
        output_s2[22]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_5_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[22]), .ZN(prince_AddKeyOut2_XORInst_5_2_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_5_3_U2 ( .A(
        prince_AddKeyOut2_XORInst_5_3_n3), .B(prince_selected_Key2_23_), .ZN(
        output_s2[23]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_5_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[23]), .ZN(prince_AddKeyOut2_XORInst_5_3_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_6_0_U2 ( .A(
        prince_AddKeyOut2_XORInst_6_0_n3), .B(prince_selected_Key2_24_), .ZN(
        output_s2[24]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_6_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[24]), .ZN(prince_AddKeyOut2_XORInst_6_0_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_6_1_U2 ( .A(
        prince_AddKeyOut2_XORInst_6_1_n3), .B(prince_selected_Key2_25_), .ZN(
        output_s2[25]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_6_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[25]), .ZN(prince_AddKeyOut2_XORInst_6_1_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_6_2_U2 ( .A(
        prince_AddKeyOut2_XORInst_6_2_n3), .B(prince_selected_Key2_26_), .ZN(
        output_s2[26]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_6_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[26]), .ZN(prince_AddKeyOut2_XORInst_6_2_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_6_3_U2 ( .A(
        prince_AddKeyOut2_XORInst_6_3_n3), .B(prince_selected_Key2_27_), .ZN(
        output_s2[27]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_6_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[27]), .ZN(prince_AddKeyOut2_XORInst_6_3_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_7_0_U2 ( .A(
        prince_AddKeyOut2_XORInst_7_0_n3), .B(prince_selected_Key2_28_), .ZN(
        output_s2[28]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_7_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[28]), .ZN(prince_AddKeyOut2_XORInst_7_0_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_7_1_U2 ( .A(
        prince_AddKeyOut2_XORInst_7_1_n3), .B(prince_selected_Key2_29_), .ZN(
        output_s2[29]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_7_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[29]), .ZN(prince_AddKeyOut2_XORInst_7_1_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_7_2_U2 ( .A(
        prince_AddKeyOut2_XORInst_7_2_n3), .B(prince_selected_Key2_30_), .ZN(
        output_s2[30]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_7_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[30]), .ZN(prince_AddKeyOut2_XORInst_7_2_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_7_3_U2 ( .A(
        prince_AddKeyOut2_XORInst_7_3_n3), .B(prince_selected_Key2_31_), .ZN(
        output_s2[31]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_7_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[31]), .ZN(prince_AddKeyOut2_XORInst_7_3_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_8_0_U2 ( .A(
        prince_AddKeyOut2_XORInst_8_0_n3), .B(prince_selected_Key2_32_), .ZN(
        output_s2[32]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_8_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[32]), .ZN(prince_AddKeyOut2_XORInst_8_0_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_8_1_U2 ( .A(
        prince_AddKeyOut2_XORInst_8_1_n3), .B(prince_selected_Key2_33_), .ZN(
        output_s2[33]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_8_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[33]), .ZN(prince_AddKeyOut2_XORInst_8_1_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_8_2_U2 ( .A(
        prince_AddKeyOut2_XORInst_8_2_n3), .B(prince_selected_Key2_34_), .ZN(
        output_s2[34]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_8_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[34]), .ZN(prince_AddKeyOut2_XORInst_8_2_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_8_3_U2 ( .A(
        prince_AddKeyOut2_XORInst_8_3_n3), .B(prince_selected_Key2_35_), .ZN(
        output_s2[35]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_8_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[35]), .ZN(prince_AddKeyOut2_XORInst_8_3_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_9_0_U2 ( .A(
        prince_AddKeyOut2_XORInst_9_0_n3), .B(prince_selected_Key2_36_), .ZN(
        output_s2[36]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_9_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[36]), .ZN(prince_AddKeyOut2_XORInst_9_0_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_9_1_U2 ( .A(
        prince_AddKeyOut2_XORInst_9_1_n3), .B(prince_selected_Key2_37_), .ZN(
        output_s2[37]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_9_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[37]), .ZN(prince_AddKeyOut2_XORInst_9_1_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_9_2_U2 ( .A(
        prince_AddKeyOut2_XORInst_9_2_n3), .B(prince_selected_Key2_38_), .ZN(
        output_s2[38]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_9_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[38]), .ZN(prince_AddKeyOut2_XORInst_9_2_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_9_3_U2 ( .A(
        prince_AddKeyOut2_XORInst_9_3_n3), .B(prince_selected_Key2_39_), .ZN(
        output_s2[39]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_9_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[39]), .ZN(prince_AddKeyOut2_XORInst_9_3_n3) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_10_0_U2 ( .A(
        prince_AddKeyOut2_XORInst_10_0_n3), .B(prince_selected_Key2_40_), .ZN(
        output_s2[40]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_10_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[40]), .ZN(prince_AddKeyOut2_XORInst_10_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_10_1_U2 ( .A(
        prince_AddKeyOut2_XORInst_10_1_n3), .B(prince_selected_Key2_41_), .ZN(
        output_s2[41]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_10_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[41]), .ZN(prince_AddKeyOut2_XORInst_10_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_10_2_U2 ( .A(
        prince_AddKeyOut2_XORInst_10_2_n3), .B(prince_selected_Key2_42_), .ZN(
        output_s2[42]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_10_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[42]), .ZN(prince_AddKeyOut2_XORInst_10_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_10_3_U2 ( .A(
        prince_AddKeyOut2_XORInst_10_3_n3), .B(prince_selected_Key2_43_), .ZN(
        output_s2[43]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_10_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[43]), .ZN(prince_AddKeyOut2_XORInst_10_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_11_0_U2 ( .A(
        prince_AddKeyOut2_XORInst_11_0_n3), .B(prince_selected_Key2_44_), .ZN(
        output_s2[44]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_11_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[44]), .ZN(prince_AddKeyOut2_XORInst_11_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_11_1_U2 ( .A(
        prince_AddKeyOut2_XORInst_11_1_n3), .B(prince_selected_Key2_45_), .ZN(
        output_s2[45]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_11_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[45]), .ZN(prince_AddKeyOut2_XORInst_11_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_11_2_U2 ( .A(
        prince_AddKeyOut2_XORInst_11_2_n3), .B(prince_selected_Key2_46_), .ZN(
        output_s2[46]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_11_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[46]), .ZN(prince_AddKeyOut2_XORInst_11_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_11_3_U2 ( .A(
        prince_AddKeyOut2_XORInst_11_3_n3), .B(prince_selected_Key2_47_), .ZN(
        output_s2[47]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_11_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[47]), .ZN(prince_AddKeyOut2_XORInst_11_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_12_0_U2 ( .A(
        prince_AddKeyOut2_XORInst_12_0_n3), .B(prince_selected_Key2_48_), .ZN(
        output_s2[48]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_12_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[48]), .ZN(prince_AddKeyOut2_XORInst_12_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_12_1_U2 ( .A(
        prince_AddKeyOut2_XORInst_12_1_n3), .B(prince_selected_Key2_49_), .ZN(
        output_s2[49]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_12_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[49]), .ZN(prince_AddKeyOut2_XORInst_12_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_12_2_U2 ( .A(
        prince_AddKeyOut2_XORInst_12_2_n3), .B(prince_selected_Key2_50_), .ZN(
        output_s2[50]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_12_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[50]), .ZN(prince_AddKeyOut2_XORInst_12_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_12_3_U2 ( .A(
        prince_AddKeyOut2_XORInst_12_3_n3), .B(prince_selected_Key2_51_), .ZN(
        output_s2[51]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_12_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[51]), .ZN(prince_AddKeyOut2_XORInst_12_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_13_0_U2 ( .A(
        prince_AddKeyOut2_XORInst_13_0_n3), .B(prince_selected_Key2_52_), .ZN(
        output_s2[52]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_13_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[52]), .ZN(prince_AddKeyOut2_XORInst_13_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_13_1_U2 ( .A(
        prince_AddKeyOut2_XORInst_13_1_n3), .B(prince_selected_Key2_53_), .ZN(
        output_s2[53]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_13_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[53]), .ZN(prince_AddKeyOut2_XORInst_13_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_13_2_U2 ( .A(
        prince_AddKeyOut2_XORInst_13_2_n3), .B(prince_selected_Key2_54_), .ZN(
        output_s2[54]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_13_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[54]), .ZN(prince_AddKeyOut2_XORInst_13_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_13_3_U2 ( .A(
        prince_AddKeyOut2_XORInst_13_3_n3), .B(prince_selected_Key2_55_), .ZN(
        output_s2[55]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_13_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[55]), .ZN(prince_AddKeyOut2_XORInst_13_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_14_0_U2 ( .A(
        prince_AddKeyOut2_XORInst_14_0_n3), .B(prince_selected_Key2_56_), .ZN(
        output_s2[56]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_14_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[56]), .ZN(prince_AddKeyOut2_XORInst_14_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_14_1_U2 ( .A(
        prince_AddKeyOut2_XORInst_14_1_n3), .B(prince_selected_Key2_57_), .ZN(
        output_s2[57]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_14_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[57]), .ZN(prince_AddKeyOut2_XORInst_14_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_14_2_U2 ( .A(
        prince_AddKeyOut2_XORInst_14_2_n3), .B(prince_selected_Key2_58_), .ZN(
        output_s2[58]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_14_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[58]), .ZN(prince_AddKeyOut2_XORInst_14_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_14_3_U2 ( .A(
        prince_AddKeyOut2_XORInst_14_3_n3), .B(prince_selected_Key2_59_), .ZN(
        output_s2[59]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_14_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[59]), .ZN(prince_AddKeyOut2_XORInst_14_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_15_0_U2 ( .A(
        prince_AddKeyOut2_XORInst_15_0_n3), .B(prince_selected_Key2_60_), .ZN(
        output_s2[60]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_15_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[60]), .ZN(prince_AddKeyOut2_XORInst_15_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_15_1_U2 ( .A(
        prince_AddKeyOut2_XORInst_15_1_n3), .B(prince_selected_Key2_61_), .ZN(
        output_s2[61]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_15_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[61]), .ZN(prince_AddKeyOut2_XORInst_15_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_15_2_U2 ( .A(
        prince_AddKeyOut2_XORInst_15_2_n3), .B(prince_selected_Key2_62_), .ZN(
        output_s2[62]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_15_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[62]), .ZN(prince_AddKeyOut2_XORInst_15_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut2_XORInst_15_3_U2 ( .A(
        prince_AddKeyOut2_XORInst_15_3_n3), .B(prince_selected_Key2_63_), .ZN(
        output_s2[63]) );
  XNOR2_X1 prince_AddKeyOut2_XORInst_15_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s2[63]), .ZN(prince_AddKeyOut2_XORInst_15_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_0_0_U2 ( .A(
        prince_AddKeyOut3_XORInst_0_0_n3), .B(prince_selected_Key3_0_), .ZN(
        output_s3[0]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_0_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[0]), .ZN(prince_AddKeyOut3_XORInst_0_0_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_0_1_U2 ( .A(
        prince_AddKeyOut3_XORInst_0_1_n3), .B(prince_selected_Key3_1_), .ZN(
        output_s3[1]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_0_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[1]), .ZN(prince_AddKeyOut3_XORInst_0_1_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_0_2_U2 ( .A(
        prince_AddKeyOut3_XORInst_0_2_n3), .B(prince_selected_Key3_2_), .ZN(
        output_s3[2]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_0_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[2]), .ZN(prince_AddKeyOut3_XORInst_0_2_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_0_3_U2 ( .A(
        prince_AddKeyOut3_XORInst_0_3_n3), .B(prince_selected_Key3_3_), .ZN(
        output_s3[3]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_0_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[3]), .ZN(prince_AddKeyOut3_XORInst_0_3_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_1_0_U2 ( .A(
        prince_AddKeyOut3_XORInst_1_0_n3), .B(prince_selected_Key3_4_), .ZN(
        output_s3[4]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_1_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[4]), .ZN(prince_AddKeyOut3_XORInst_1_0_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_1_1_U2 ( .A(
        prince_AddKeyOut3_XORInst_1_1_n3), .B(prince_selected_Key3_5_), .ZN(
        output_s3[5]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_1_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[5]), .ZN(prince_AddKeyOut3_XORInst_1_1_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_1_2_U2 ( .A(
        prince_AddKeyOut3_XORInst_1_2_n3), .B(prince_selected_Key3_6_), .ZN(
        output_s3[6]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_1_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[6]), .ZN(prince_AddKeyOut3_XORInst_1_2_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_1_3_U2 ( .A(
        prince_AddKeyOut3_XORInst_1_3_n3), .B(prince_selected_Key3_7_), .ZN(
        output_s3[7]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_1_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[7]), .ZN(prince_AddKeyOut3_XORInst_1_3_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_2_0_U2 ( .A(
        prince_AddKeyOut3_XORInst_2_0_n3), .B(prince_selected_Key3_8_), .ZN(
        output_s3[8]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_2_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[8]), .ZN(prince_AddKeyOut3_XORInst_2_0_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_2_1_U2 ( .A(
        prince_AddKeyOut3_XORInst_2_1_n3), .B(prince_selected_Key3_9_), .ZN(
        output_s3[9]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_2_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[9]), .ZN(prince_AddKeyOut3_XORInst_2_1_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_2_2_U2 ( .A(
        prince_AddKeyOut3_XORInst_2_2_n3), .B(prince_selected_Key3_10_), .ZN(
        output_s3[10]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_2_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[10]), .ZN(prince_AddKeyOut3_XORInst_2_2_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_2_3_U2 ( .A(
        prince_AddKeyOut3_XORInst_2_3_n3), .B(prince_selected_Key3_11_), .ZN(
        output_s3[11]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_2_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[11]), .ZN(prince_AddKeyOut3_XORInst_2_3_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_3_0_U2 ( .A(
        prince_AddKeyOut3_XORInst_3_0_n3), .B(prince_selected_Key3_12_), .ZN(
        output_s3[12]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_3_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[12]), .ZN(prince_AddKeyOut3_XORInst_3_0_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_3_1_U2 ( .A(
        prince_AddKeyOut3_XORInst_3_1_n3), .B(prince_selected_Key3_13_), .ZN(
        output_s3[13]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_3_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[13]), .ZN(prince_AddKeyOut3_XORInst_3_1_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_3_2_U2 ( .A(
        prince_AddKeyOut3_XORInst_3_2_n3), .B(prince_selected_Key3_14_), .ZN(
        output_s3[14]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_3_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[14]), .ZN(prince_AddKeyOut3_XORInst_3_2_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_3_3_U2 ( .A(
        prince_AddKeyOut3_XORInst_3_3_n3), .B(prince_selected_Key3_15_), .ZN(
        output_s3[15]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_3_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[15]), .ZN(prince_AddKeyOut3_XORInst_3_3_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_4_0_U2 ( .A(
        prince_AddKeyOut3_XORInst_4_0_n3), .B(prince_selected_Key3_16_), .ZN(
        output_s3[16]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_4_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[16]), .ZN(prince_AddKeyOut3_XORInst_4_0_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_4_1_U2 ( .A(
        prince_AddKeyOut3_XORInst_4_1_n3), .B(prince_selected_Key3_17_), .ZN(
        output_s3[17]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_4_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[17]), .ZN(prince_AddKeyOut3_XORInst_4_1_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_4_2_U2 ( .A(
        prince_AddKeyOut3_XORInst_4_2_n3), .B(prince_selected_Key3_18_), .ZN(
        output_s3[18]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_4_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[18]), .ZN(prince_AddKeyOut3_XORInst_4_2_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_4_3_U2 ( .A(
        prince_AddKeyOut3_XORInst_4_3_n3), .B(prince_selected_Key3_19_), .ZN(
        output_s3[19]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_4_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[19]), .ZN(prince_AddKeyOut3_XORInst_4_3_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_5_0_U2 ( .A(
        prince_AddKeyOut3_XORInst_5_0_n3), .B(prince_selected_Key3_20_), .ZN(
        output_s3[20]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_5_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[20]), .ZN(prince_AddKeyOut3_XORInst_5_0_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_5_1_U2 ( .A(
        prince_AddKeyOut3_XORInst_5_1_n3), .B(prince_selected_Key3_21_), .ZN(
        output_s3[21]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_5_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[21]), .ZN(prince_AddKeyOut3_XORInst_5_1_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_5_2_U2 ( .A(
        prince_AddKeyOut3_XORInst_5_2_n3), .B(prince_selected_Key3_22_), .ZN(
        output_s3[22]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_5_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[22]), .ZN(prince_AddKeyOut3_XORInst_5_2_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_5_3_U2 ( .A(
        prince_AddKeyOut3_XORInst_5_3_n3), .B(prince_selected_Key3_23_), .ZN(
        output_s3[23]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_5_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[23]), .ZN(prince_AddKeyOut3_XORInst_5_3_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_6_0_U2 ( .A(
        prince_AddKeyOut3_XORInst_6_0_n3), .B(prince_selected_Key3_24_), .ZN(
        output_s3[24]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_6_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[24]), .ZN(prince_AddKeyOut3_XORInst_6_0_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_6_1_U2 ( .A(
        prince_AddKeyOut3_XORInst_6_1_n3), .B(prince_selected_Key3_25_), .ZN(
        output_s3[25]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_6_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[25]), .ZN(prince_AddKeyOut3_XORInst_6_1_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_6_2_U2 ( .A(
        prince_AddKeyOut3_XORInst_6_2_n3), .B(prince_selected_Key3_26_), .ZN(
        output_s3[26]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_6_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[26]), .ZN(prince_AddKeyOut3_XORInst_6_2_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_6_3_U2 ( .A(
        prince_AddKeyOut3_XORInst_6_3_n3), .B(prince_selected_Key3_27_), .ZN(
        output_s3[27]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_6_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[27]), .ZN(prince_AddKeyOut3_XORInst_6_3_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_7_0_U2 ( .A(
        prince_AddKeyOut3_XORInst_7_0_n3), .B(prince_selected_Key3_28_), .ZN(
        output_s3[28]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_7_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[28]), .ZN(prince_AddKeyOut3_XORInst_7_0_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_7_1_U2 ( .A(
        prince_AddKeyOut3_XORInst_7_1_n3), .B(prince_selected_Key3_29_), .ZN(
        output_s3[29]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_7_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[29]), .ZN(prince_AddKeyOut3_XORInst_7_1_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_7_2_U2 ( .A(
        prince_AddKeyOut3_XORInst_7_2_n3), .B(prince_selected_Key3_30_), .ZN(
        output_s3[30]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_7_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[30]), .ZN(prince_AddKeyOut3_XORInst_7_2_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_7_3_U2 ( .A(
        prince_AddKeyOut3_XORInst_7_3_n3), .B(prince_selected_Key3_31_), .ZN(
        output_s3[31]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_7_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[31]), .ZN(prince_AddKeyOut3_XORInst_7_3_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_8_0_U2 ( .A(
        prince_AddKeyOut3_XORInst_8_0_n3), .B(prince_selected_Key3_32_), .ZN(
        output_s3[32]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_8_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[32]), .ZN(prince_AddKeyOut3_XORInst_8_0_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_8_1_U2 ( .A(
        prince_AddKeyOut3_XORInst_8_1_n3), .B(prince_selected_Key3_33_), .ZN(
        output_s3[33]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_8_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[33]), .ZN(prince_AddKeyOut3_XORInst_8_1_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_8_2_U2 ( .A(
        prince_AddKeyOut3_XORInst_8_2_n3), .B(prince_selected_Key3_34_), .ZN(
        output_s3[34]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_8_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[34]), .ZN(prince_AddKeyOut3_XORInst_8_2_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_8_3_U2 ( .A(
        prince_AddKeyOut3_XORInst_8_3_n3), .B(prince_selected_Key3_35_), .ZN(
        output_s3[35]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_8_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[35]), .ZN(prince_AddKeyOut3_XORInst_8_3_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_9_0_U2 ( .A(
        prince_AddKeyOut3_XORInst_9_0_n3), .B(prince_selected_Key3_36_), .ZN(
        output_s3[36]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_9_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[36]), .ZN(prince_AddKeyOut3_XORInst_9_0_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_9_1_U2 ( .A(
        prince_AddKeyOut3_XORInst_9_1_n3), .B(prince_selected_Key3_37_), .ZN(
        output_s3[37]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_9_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[37]), .ZN(prince_AddKeyOut3_XORInst_9_1_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_9_2_U2 ( .A(
        prince_AddKeyOut3_XORInst_9_2_n3), .B(prince_selected_Key3_38_), .ZN(
        output_s3[38]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_9_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[38]), .ZN(prince_AddKeyOut3_XORInst_9_2_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_9_3_U2 ( .A(
        prince_AddKeyOut3_XORInst_9_3_n3), .B(prince_selected_Key3_39_), .ZN(
        output_s3[39]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_9_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[39]), .ZN(prince_AddKeyOut3_XORInst_9_3_n3) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_10_0_U2 ( .A(
        prince_AddKeyOut3_XORInst_10_0_n3), .B(prince_selected_Key3_40_), .ZN(
        output_s3[40]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_10_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[40]), .ZN(prince_AddKeyOut3_XORInst_10_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_10_1_U2 ( .A(
        prince_AddKeyOut3_XORInst_10_1_n3), .B(prince_selected_Key3_41_), .ZN(
        output_s3[41]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_10_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[41]), .ZN(prince_AddKeyOut3_XORInst_10_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_10_2_U2 ( .A(
        prince_AddKeyOut3_XORInst_10_2_n3), .B(prince_selected_Key3_42_), .ZN(
        output_s3[42]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_10_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[42]), .ZN(prince_AddKeyOut3_XORInst_10_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_10_3_U2 ( .A(
        prince_AddKeyOut3_XORInst_10_3_n3), .B(prince_selected_Key3_43_), .ZN(
        output_s3[43]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_10_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[43]), .ZN(prince_AddKeyOut3_XORInst_10_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_11_0_U2 ( .A(
        prince_AddKeyOut3_XORInst_11_0_n3), .B(prince_selected_Key3_44_), .ZN(
        output_s3[44]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_11_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[44]), .ZN(prince_AddKeyOut3_XORInst_11_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_11_1_U2 ( .A(
        prince_AddKeyOut3_XORInst_11_1_n3), .B(prince_selected_Key3_45_), .ZN(
        output_s3[45]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_11_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[45]), .ZN(prince_AddKeyOut3_XORInst_11_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_11_2_U2 ( .A(
        prince_AddKeyOut3_XORInst_11_2_n3), .B(prince_selected_Key3_46_), .ZN(
        output_s3[46]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_11_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[46]), .ZN(prince_AddKeyOut3_XORInst_11_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_11_3_U2 ( .A(
        prince_AddKeyOut3_XORInst_11_3_n3), .B(prince_selected_Key3_47_), .ZN(
        output_s3[47]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_11_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[47]), .ZN(prince_AddKeyOut3_XORInst_11_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_12_0_U2 ( .A(
        prince_AddKeyOut3_XORInst_12_0_n3), .B(prince_selected_Key3_48_), .ZN(
        output_s3[48]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_12_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[48]), .ZN(prince_AddKeyOut3_XORInst_12_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_12_1_U2 ( .A(
        prince_AddKeyOut3_XORInst_12_1_n3), .B(prince_selected_Key3_49_), .ZN(
        output_s3[49]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_12_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[49]), .ZN(prince_AddKeyOut3_XORInst_12_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_12_2_U2 ( .A(
        prince_AddKeyOut3_XORInst_12_2_n3), .B(prince_selected_Key3_50_), .ZN(
        output_s3[50]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_12_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[50]), .ZN(prince_AddKeyOut3_XORInst_12_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_12_3_U2 ( .A(
        prince_AddKeyOut3_XORInst_12_3_n3), .B(prince_selected_Key3_51_), .ZN(
        output_s3[51]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_12_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[51]), .ZN(prince_AddKeyOut3_XORInst_12_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_13_0_U2 ( .A(
        prince_AddKeyOut3_XORInst_13_0_n3), .B(prince_selected_Key3_52_), .ZN(
        output_s3[52]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_13_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[52]), .ZN(prince_AddKeyOut3_XORInst_13_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_13_1_U2 ( .A(
        prince_AddKeyOut3_XORInst_13_1_n3), .B(prince_selected_Key3_53_), .ZN(
        output_s3[53]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_13_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[53]), .ZN(prince_AddKeyOut3_XORInst_13_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_13_2_U2 ( .A(
        prince_AddKeyOut3_XORInst_13_2_n3), .B(prince_selected_Key3_54_), .ZN(
        output_s3[54]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_13_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[54]), .ZN(prince_AddKeyOut3_XORInst_13_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_13_3_U2 ( .A(
        prince_AddKeyOut3_XORInst_13_3_n3), .B(prince_selected_Key3_55_), .ZN(
        output_s3[55]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_13_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[55]), .ZN(prince_AddKeyOut3_XORInst_13_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_14_0_U2 ( .A(
        prince_AddKeyOut3_XORInst_14_0_n3), .B(prince_selected_Key3_56_), .ZN(
        output_s3[56]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_14_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[56]), .ZN(prince_AddKeyOut3_XORInst_14_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_14_1_U2 ( .A(
        prince_AddKeyOut3_XORInst_14_1_n3), .B(prince_selected_Key3_57_), .ZN(
        output_s3[57]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_14_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[57]), .ZN(prince_AddKeyOut3_XORInst_14_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_14_2_U2 ( .A(
        prince_AddKeyOut3_XORInst_14_2_n3), .B(prince_selected_Key3_58_), .ZN(
        output_s3[58]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_14_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[58]), .ZN(prince_AddKeyOut3_XORInst_14_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_14_3_U2 ( .A(
        prince_AddKeyOut3_XORInst_14_3_n3), .B(prince_selected_Key3_59_), .ZN(
        output_s3[59]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_14_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[59]), .ZN(prince_AddKeyOut3_XORInst_14_3_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_15_0_U2 ( .A(
        prince_AddKeyOut3_XORInst_15_0_n3), .B(prince_selected_Key3_60_), .ZN(
        output_s3[60]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_15_0_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[60]), .ZN(prince_AddKeyOut3_XORInst_15_0_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_15_1_U2 ( .A(
        prince_AddKeyOut3_XORInst_15_1_n3), .B(prince_selected_Key3_61_), .ZN(
        output_s3[61]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_15_1_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[61]), .ZN(prince_AddKeyOut3_XORInst_15_1_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_15_2_U2 ( .A(
        prince_AddKeyOut3_XORInst_15_2_n3), .B(prince_selected_Key3_62_), .ZN(
        output_s3[62]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_15_2_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[62]), .ZN(prince_AddKeyOut3_XORInst_15_2_n3)
         );
  XNOR2_X1 prince_AddKeyOut3_XORInst_15_3_U2 ( .A(
        prince_AddKeyOut3_XORInst_15_3_n3), .B(prince_selected_Key3_63_), .ZN(
        output_s3[63]) );
  XNOR2_X1 prince_AddKeyOut3_XORInst_15_3_U1 ( .A(1'b0), .B(
        prince_rounds_Output_s3[63]), .ZN(prince_AddKeyOut3_XORInst_15_3_n3)
         );
endmodule

