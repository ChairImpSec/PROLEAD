module circuit ( sboxIn, randomS2, randomS3, randomS4, randomS5, clk, sboxOut );
  input [15:0] sboxIn;
  input [15:0] randomS2;
  input [7:0] randomS3;
  input [15:0] randomS4;
  input [31:0] randomS5;
  output [15:0] sboxOut;
  input clk;
  wire   s1_linMapOut_0__0_, s1_linMapOut_0__1_, s1_linMapOut_0__3_,
         s1_linMapOut_0__4_, s1_linMapOut_0__5_, s1_linMapOut_0__6_,
         s1_linMapOut_0__7_, s1_linMapOut_1__0_, s1_linMapOut_1__1_,
         s1_linMapOut_1__3_, s1_linMapOut_1__4_, s1_linMapOut_1__5_,
         s1_linMapOut_1__6_, s1_linMapOut_1__7_, s1_input_mapping_1_n23,
         s1_input_mapping_1_n22, s1_input_mapping_1_n21,
         s1_input_mapping_1_n20, s1_input_mapping_1_n19,
         s1_input_mapping_1_n18, s1_input_mapping_1_n17,
         s1_input_mapping_0_n23, s1_input_mapping_0_n22,
         s1_input_mapping_0_n21, s1_input_mapping_0_n20,
         s1_input_mapping_0_n19, s1_input_mapping_0_n18,
         s1_input_mapping_0_n17, s2_n16, s2_n15, s2_n14, s2_n13, s2_n12,
         s2_n11, s2_n10, s2_n9, s2_n8, s2_n7, s2_n6, s2_n5, s2_n4, s2_n3,
         s2_n2, s2_n1, s2_regOut_0__1__0_, s2_regOut_0__1__1_,
         s2_regOut_0__1__2_, s2_regOut_0__1__3_, s2_regOut_0__2__0_,
         s2_regOut_0__2__1_, s2_regOut_0__2__2_, s2_regOut_0__2__3_,
         s2_regOut_1__1__0_, s2_regOut_1__1__1_, s2_regOut_1__1__2_,
         s2_regOut_1__1__3_, s2_regOut_1__2__0_, s2_regOut_1__2__1_,
         s2_regOut_1__2__2_, s2_regOut_1__2__3_, s2_gf2_mul_out_0__0__0_,
         s2_gf2_mul_out_0__0__1_, s2_gf2_mul_out_0__0__2_,
         s2_gf2_mul_out_0__0__3_, s2_gf2_mul_out_1__1__0_,
         s2_gf2_mul_out_1__1__1_, s2_gf2_mul_out_1__1__2_,
         s2_gf2_mul_out_1__1__3_, s2_sqsc_in_0__0_, s2_sqsc_in_0__1_,
         s2_sqsc_in_0__2_, s2_sqsc_in_0__3_, s2_sqsc_in_1__0_,
         s2_sqsc_in_1__1_, s2_sqsc_in_1__2_, s2_sqsc_in_1__3_, s2_mul1_1_1_n77,
         s2_mul1_1_1_n76, s2_mul1_1_1_n75, s2_mul1_1_1_n74, s2_mul1_1_1_n73,
         s2_mul1_1_1_n72, s2_mul1_1_1_n71, s2_mul1_1_1_n70, s2_mul1_1_1_n69,
         s2_mul1_1_1_n68, s2_mul1_1_1_n67, s2_mul1_1_1_n66, s2_mul1_1_1_n65,
         s2_mul1_1_1_n64, s2_mul1_1_1_n63, s2_mul1_1_1_n62, s2_mul1_1_1_n61,
         s2_mul1_1_1_n60, s2_mul1_1_1_n59, s2_mul1_1_1_n58, s2_mul1_1_1_n57,
         s2_mul1_1_1_n56, s2_mul1_1_1_n55, s2_mul1_1_1_n54, s2_mul1_1_1_n53,
         s2_mul1_1_0_n77, s2_mul1_1_0_n76, s2_mul1_1_0_n75, s2_mul1_1_0_n74,
         s2_mul1_1_0_n73, s2_mul1_1_0_n72, s2_mul1_1_0_n71, s2_mul1_1_0_n70,
         s2_mul1_1_0_n69, s2_mul1_1_0_n68, s2_mul1_1_0_n67, s2_mul1_1_0_n66,
         s2_mul1_1_0_n65, s2_mul1_1_0_n64, s2_mul1_1_0_n63, s2_mul1_1_0_n62,
         s2_mul1_1_0_n61, s2_mul1_1_0_n60, s2_mul1_1_0_n59, s2_mul1_1_0_n58,
         s2_mul1_1_0_n57, s2_mul1_1_0_n56, s2_mul1_1_0_n55, s2_mul1_1_0_n54,
         s2_mul1_1_0_n53, s2_mul1_0_1_n77, s2_mul1_0_1_n76, s2_mul1_0_1_n75,
         s2_mul1_0_1_n74, s2_mul1_0_1_n73, s2_mul1_0_1_n72, s2_mul1_0_1_n71,
         s2_mul1_0_1_n70, s2_mul1_0_1_n69, s2_mul1_0_1_n68, s2_mul1_0_1_n67,
         s2_mul1_0_1_n66, s2_mul1_0_1_n65, s2_mul1_0_1_n64, s2_mul1_0_1_n63,
         s2_mul1_0_1_n62, s2_mul1_0_1_n61, s2_mul1_0_1_n60, s2_mul1_0_1_n59,
         s2_mul1_0_1_n58, s2_mul1_0_1_n57, s2_mul1_0_1_n56, s2_mul1_0_1_n55,
         s2_mul1_0_1_n54, s2_mul1_0_1_n53, s2_mul1_0_0_n77, s2_mul1_0_0_n76,
         s2_mul1_0_0_n75, s2_mul1_0_0_n74, s2_mul1_0_0_n73, s2_mul1_0_0_n72,
         s2_mul1_0_0_n71, s2_mul1_0_0_n70, s2_mul1_0_0_n69, s2_mul1_0_0_n68,
         s2_mul1_0_0_n67, s2_mul1_0_0_n66, s2_mul1_0_0_n65, s2_mul1_0_0_n64,
         s2_mul1_0_0_n63, s2_mul1_0_0_n62, s2_mul1_0_0_n61, s2_mul1_0_0_n60,
         s2_mul1_0_0_n59, s2_mul1_0_0_n58, s2_mul1_0_0_n57, s2_mul1_0_0_n56,
         s2_mul1_0_0_n55, s2_mul1_0_0_n54, s2_mul1_0_0_n53, s3_n8, s3_n7,
         s3_n6, s3_n5, s3_n4, s3_n3, s3_n2, s3_n1, s3_regOut_0__3__0_,
         s3_regOut_0__3__1_, s3_regOut_0__4__0_, s3_regOut_0__4__1_,
         s3_regOut_1__3__0_, s3_regOut_1__3__1_, s3_regOut_1__4__0_,
         s3_regOut_1__4__1_, s3_gf2_mul_out_0__0__0_, s3_gf2_mul_out_0__0__1_,
         s3_gf2_mul_out_1__1__0_, s3_gf2_mul_out_1__1__1_, s3_scale_in_0__0_,
         s3_scale_in_0__1_, s3_scale_in_1__0_, s3_scale_in_1__1_,
         s3_mul1_1_1_n15, s3_mul1_1_1_n14, s3_mul1_1_1_n13, s3_mul1_1_1_n12,
         s3_mul1_1_1_n11, s3_mul1_1_0_n15, s3_mul1_1_0_n14, s3_mul1_1_0_n13,
         s3_mul1_1_0_n12, s3_mul1_1_0_n11, s3_mul1_0_1_n15, s3_mul1_0_1_n14,
         s3_mul1_0_1_n13, s3_mul1_0_1_n12, s3_mul1_0_1_n11, s3_mul1_0_0_n15,
         s3_mul1_0_0_n14, s3_mul1_0_0_n13, s3_mul1_0_0_n12, s3_mul1_0_0_n11,
         s4_n8, s4_n7, s4_n6, s4_n5, s4_n4, s4_n3, s4_n2, s4_n1,
         s4_regOut_0__1__0_, s4_regOut_0__1__1_, s4_regOut_0__1__2_,
         s4_regOut_0__1__3_, s4_regOut_0__2__0_, s4_regOut_0__2__1_,
         s4_regOut_0__2__2_, s4_regOut_0__2__3_, s4_regOut_1__1__0_,
         s4_regOut_1__1__1_, s4_regOut_1__1__2_, s4_regOut_1__1__3_,
         s4_regOut_1__2__0_, s4_regOut_1__2__1_, s4_regOut_1__2__2_,
         s4_regOut_1__2__3_, s4_inv_out_0__0_, s4_inv_out_0__1_,
         s4_inv_out_1__0_, s4_inv_out_1__1_, s4_mul1_1_1_n15, s4_mul1_1_1_n14,
         s4_mul1_1_1_n13, s4_mul1_1_1_n12, s4_mul1_1_1_n11, s4_mul1_1_0_n15,
         s4_mul1_1_0_n14, s4_mul1_1_0_n13, s4_mul1_1_0_n12, s4_mul1_1_0_n11,
         s4_mul1_0_1_n15, s4_mul1_0_1_n14, s4_mul1_0_1_n13, s4_mul1_0_1_n12,
         s4_mul1_0_1_n11, s4_mul1_0_0_n15, s4_mul1_0_0_n14, s4_mul1_0_0_n13,
         s4_mul1_0_0_n12, s4_mul1_0_0_n11, s4_mul2_1_1_n15, s4_mul2_1_1_n14,
         s4_mul2_1_1_n13, s4_mul2_1_1_n12, s4_mul2_1_1_n11, s4_mul2_1_0_n15,
         s4_mul2_1_0_n14, s4_mul2_1_0_n13, s4_mul2_1_0_n12, s4_mul2_1_0_n11,
         s4_mul2_0_1_n15, s4_mul2_0_1_n14, s4_mul2_0_1_n13, s4_mul2_0_1_n12,
         s4_mul2_0_1_n11, s4_mul2_0_0_n15, s4_mul2_0_0_n14, s4_mul2_0_0_n13,
         s4_mul2_0_0_n12, s4_mul2_0_0_n11, s5_n16, s5_n15, s5_n14, s5_n13,
         s5_n12, s5_n11, s5_n10, s5_n9, s5_n8, s5_n7, s5_n6, s5_n5, s5_n4,
         s5_n3, s5_n2, s5_n1, s5_mul1_1_1_n77, s5_mul1_1_1_n76,
         s5_mul1_1_1_n75, s5_mul1_1_1_n74, s5_mul1_1_1_n73, s5_mul1_1_1_n72,
         s5_mul1_1_1_n71, s5_mul1_1_1_n70, s5_mul1_1_1_n69, s5_mul1_1_1_n68,
         s5_mul1_1_1_n67, s5_mul1_1_1_n66, s5_mul1_1_1_n65, s5_mul1_1_1_n64,
         s5_mul1_1_1_n63, s5_mul1_1_1_n62, s5_mul1_1_1_n61, s5_mul1_1_1_n60,
         s5_mul1_1_1_n59, s5_mul1_1_1_n58, s5_mul1_1_1_n57, s5_mul1_1_1_n56,
         s5_mul1_1_1_n55, s5_mul1_1_1_n54, s5_mul1_1_1_n53, s5_mul1_1_0_n77,
         s5_mul1_1_0_n76, s5_mul1_1_0_n75, s5_mul1_1_0_n74, s5_mul1_1_0_n73,
         s5_mul1_1_0_n72, s5_mul1_1_0_n71, s5_mul1_1_0_n70, s5_mul1_1_0_n69,
         s5_mul1_1_0_n68, s5_mul1_1_0_n67, s5_mul1_1_0_n66, s5_mul1_1_0_n65,
         s5_mul1_1_0_n64, s5_mul1_1_0_n63, s5_mul1_1_0_n62, s5_mul1_1_0_n61,
         s5_mul1_1_0_n60, s5_mul1_1_0_n59, s5_mul1_1_0_n58, s5_mul1_1_0_n57,
         s5_mul1_1_0_n56, s5_mul1_1_0_n55, s5_mul1_1_0_n54, s5_mul1_1_0_n53,
         s5_mul1_0_1_n77, s5_mul1_0_1_n76, s5_mul1_0_1_n75, s5_mul1_0_1_n74,
         s5_mul1_0_1_n73, s5_mul1_0_1_n72, s5_mul1_0_1_n71, s5_mul1_0_1_n70,
         s5_mul1_0_1_n69, s5_mul1_0_1_n68, s5_mul1_0_1_n67, s5_mul1_0_1_n66,
         s5_mul1_0_1_n65, s5_mul1_0_1_n64, s5_mul1_0_1_n63, s5_mul1_0_1_n62,
         s5_mul1_0_1_n61, s5_mul1_0_1_n60, s5_mul1_0_1_n59, s5_mul1_0_1_n58,
         s5_mul1_0_1_n57, s5_mul1_0_1_n56, s5_mul1_0_1_n55, s5_mul1_0_1_n54,
         s5_mul1_0_1_n53, s5_mul1_0_0_n77, s5_mul1_0_0_n76, s5_mul1_0_0_n75,
         s5_mul1_0_0_n74, s5_mul1_0_0_n73, s5_mul1_0_0_n72, s5_mul1_0_0_n71,
         s5_mul1_0_0_n70, s5_mul1_0_0_n69, s5_mul1_0_0_n68, s5_mul1_0_0_n67,
         s5_mul1_0_0_n66, s5_mul1_0_0_n65, s5_mul1_0_0_n64, s5_mul1_0_0_n63,
         s5_mul1_0_0_n62, s5_mul1_0_0_n61, s5_mul1_0_0_n60, s5_mul1_0_0_n59,
         s5_mul1_0_0_n58, s5_mul1_0_0_n57, s5_mul1_0_0_n56, s5_mul1_0_0_n55,
         s5_mul1_0_0_n54, s5_mul1_0_0_n53, s5_mul2_1_1_n77, s5_mul2_1_1_n76,
         s5_mul2_1_1_n75, s5_mul2_1_1_n74, s5_mul2_1_1_n73, s5_mul2_1_1_n72,
         s5_mul2_1_1_n71, s5_mul2_1_1_n70, s5_mul2_1_1_n69, s5_mul2_1_1_n68,
         s5_mul2_1_1_n67, s5_mul2_1_1_n66, s5_mul2_1_1_n65, s5_mul2_1_1_n64,
         s5_mul2_1_1_n63, s5_mul2_1_1_n62, s5_mul2_1_1_n61, s5_mul2_1_1_n60,
         s5_mul2_1_1_n59, s5_mul2_1_1_n58, s5_mul2_1_1_n57, s5_mul2_1_1_n56,
         s5_mul2_1_1_n55, s5_mul2_1_1_n54, s5_mul2_1_1_n53, s5_mul2_1_0_n77,
         s5_mul2_1_0_n76, s5_mul2_1_0_n75, s5_mul2_1_0_n74, s5_mul2_1_0_n73,
         s5_mul2_1_0_n72, s5_mul2_1_0_n71, s5_mul2_1_0_n70, s5_mul2_1_0_n69,
         s5_mul2_1_0_n68, s5_mul2_1_0_n67, s5_mul2_1_0_n66, s5_mul2_1_0_n65,
         s5_mul2_1_0_n64, s5_mul2_1_0_n63, s5_mul2_1_0_n62, s5_mul2_1_0_n61,
         s5_mul2_1_0_n60, s5_mul2_1_0_n59, s5_mul2_1_0_n58, s5_mul2_1_0_n57,
         s5_mul2_1_0_n56, s5_mul2_1_0_n55, s5_mul2_1_0_n54, s5_mul2_1_0_n53,
         s5_mul2_0_1_n77, s5_mul2_0_1_n76, s5_mul2_0_1_n75, s5_mul2_0_1_n74,
         s5_mul2_0_1_n73, s5_mul2_0_1_n72, s5_mul2_0_1_n71, s5_mul2_0_1_n70,
         s5_mul2_0_1_n69, s5_mul2_0_1_n68, s5_mul2_0_1_n67, s5_mul2_0_1_n66,
         s5_mul2_0_1_n65, s5_mul2_0_1_n64, s5_mul2_0_1_n63, s5_mul2_0_1_n62,
         s5_mul2_0_1_n61, s5_mul2_0_1_n60, s5_mul2_0_1_n59, s5_mul2_0_1_n58,
         s5_mul2_0_1_n57, s5_mul2_0_1_n56, s5_mul2_0_1_n55, s5_mul2_0_1_n54,
         s5_mul2_0_1_n53, s5_mul2_0_0_n77, s5_mul2_0_0_n76, s5_mul2_0_0_n75,
         s5_mul2_0_0_n74, s5_mul2_0_0_n73, s5_mul2_0_0_n72, s5_mul2_0_0_n71,
         s5_mul2_0_0_n70, s5_mul2_0_0_n69, s5_mul2_0_0_n68, s5_mul2_0_0_n67,
         s5_mul2_0_0_n66, s5_mul2_0_0_n65, s5_mul2_0_0_n64, s5_mul2_0_0_n63,
         s5_mul2_0_0_n62, s5_mul2_0_0_n61, s5_mul2_0_0_n60, s5_mul2_0_0_n59,
         s5_mul2_0_0_n58, s5_mul2_0_0_n57, s5_mul2_0_0_n56, s5_mul2_0_0_n55,
         s5_mul2_0_0_n54, s5_mul2_0_0_n53, s6_1_n9, s6_1_n8, s6_1_n7, s6_0_n9,
         s6_0_n8, s6_0_n7;
  wire   [15:0] stage1Out;
  wire   [23:0] stage2Out;
  wire   [23:0] stage3Out;
  wire   [23:0] stage4Out;
  wire   [15:0] stage5Out;
  wire   [15:0] stage6Out;
  wire   [15:0] regOut1;
  wire   [15:0] s2_refreshed;
  wire   [7:0] s2_xorResult;
  wire   [5:0] s2_sqsc_out;
  wire   [7:0] s3_refreshed;
  wire   [3:0] s3_xorResult;
  wire   [1:0] s3_scale_out;
  wire   [15:0] s4_refreshed;
  wire   [15:0] s4_concat;
  wire   [31:0] s5_regOut;
  wire   [31:0] s5_refreshed;
  wire   [31:0] s5_concat;

  DFF_X1 regOut1_reg_1__7_ ( .D(stage6Out[15]), .CK(clk), .Q(regOut1[15]), 
        .QN() );
  DFF_X1 regOut2_reg_1__7_ ( .D(regOut1[15]), .CK(clk), .Q(sboxOut[15]), .QN()
         );
  DFF_X1 regOut1_reg_1__6_ ( .D(stage6Out[14]), .CK(clk), .Q(regOut1[14]), 
        .QN() );
  DFF_X1 regOut2_reg_1__6_ ( .D(regOut1[14]), .CK(clk), .Q(sboxOut[14]), .QN()
         );
  DFF_X1 regOut1_reg_1__5_ ( .D(stage6Out[13]), .CK(clk), .Q(regOut1[13]), 
        .QN() );
  DFF_X1 regOut2_reg_1__5_ ( .D(regOut1[13]), .CK(clk), .Q(sboxOut[13]), .QN()
         );
  DFF_X1 regOut1_reg_1__4_ ( .D(stage6Out[12]), .CK(clk), .Q(regOut1[12]), 
        .QN() );
  DFF_X1 regOut2_reg_1__4_ ( .D(regOut1[12]), .CK(clk), .Q(sboxOut[12]), .QN()
         );
  DFF_X1 regOut1_reg_1__3_ ( .D(stage6Out[11]), .CK(clk), .Q(regOut1[11]), 
        .QN() );
  DFF_X1 regOut2_reg_1__3_ ( .D(regOut1[11]), .CK(clk), .Q(sboxOut[11]), .QN()
         );
  DFF_X1 regOut1_reg_1__2_ ( .D(stage6Out[10]), .CK(clk), .Q(regOut1[10]), 
        .QN() );
  DFF_X1 regOut2_reg_1__2_ ( .D(regOut1[10]), .CK(clk), .Q(sboxOut[10]), .QN()
         );
  DFF_X1 regOut1_reg_1__1_ ( .D(stage6Out[9]), .CK(clk), .Q(regOut1[9]), .QN()
         );
  DFF_X1 regOut2_reg_1__1_ ( .D(regOut1[9]), .CK(clk), .Q(sboxOut[9]), .QN()
         );
  DFF_X1 regOut1_reg_1__0_ ( .D(stage6Out[8]), .CK(clk), .Q(regOut1[8]), .QN()
         );
  DFF_X1 regOut2_reg_1__0_ ( .D(regOut1[8]), .CK(clk), .Q(sboxOut[8]), .QN()
         );
  DFF_X1 regOut1_reg_0__7_ ( .D(stage6Out[7]), .CK(clk), .Q(regOut1[7]), .QN()
         );
  DFF_X1 regOut2_reg_0__7_ ( .D(regOut1[7]), .CK(clk), .Q(sboxOut[7]), .QN()
         );
  DFF_X1 regOut1_reg_0__6_ ( .D(stage6Out[6]), .CK(clk), .Q(regOut1[6]), .QN()
         );
  DFF_X1 regOut2_reg_0__6_ ( .D(regOut1[6]), .CK(clk), .Q(), .QN(sboxOut[6])
         );
  DFF_X1 regOut1_reg_0__5_ ( .D(stage6Out[5]), .CK(clk), .Q(regOut1[5]), .QN()
         );
  DFF_X1 regOut2_reg_0__5_ ( .D(regOut1[5]), .CK(clk), .Q(), .QN(sboxOut[5])
         );
  DFF_X1 regOut1_reg_0__4_ ( .D(stage6Out[4]), .CK(clk), .Q(regOut1[4]), .QN()
         );
  DFF_X1 regOut2_reg_0__4_ ( .D(regOut1[4]), .CK(clk), .Q(sboxOut[4]), .QN()
         );
  DFF_X1 regOut1_reg_0__3_ ( .D(stage6Out[3]), .CK(clk), .Q(regOut1[3]), .QN()
         );
  DFF_X1 regOut2_reg_0__3_ ( .D(regOut1[3]), .CK(clk), .Q(sboxOut[3]), .QN()
         );
  DFF_X1 regOut1_reg_0__2_ ( .D(stage6Out[2]), .CK(clk), .Q(regOut1[2]), .QN()
         );
  DFF_X1 regOut2_reg_0__2_ ( .D(regOut1[2]), .CK(clk), .Q(sboxOut[2]), .QN()
         );
  DFF_X1 regOut1_reg_0__1_ ( .D(stage6Out[1]), .CK(clk), .Q(regOut1[1]), .QN()
         );
  DFF_X1 regOut2_reg_0__1_ ( .D(regOut1[1]), .CK(clk), .Q(), .QN(sboxOut[1])
         );
  DFF_X1 regOut1_reg_0__0_ ( .D(stage6Out[0]), .CK(clk), .Q(regOut1[0]), .QN()
         );
  DFF_X1 regOut2_reg_0__0_ ( .D(regOut1[0]), .CK(clk), .Q(), .QN(sboxOut[0])
         );
  DFF_X1 s1_stage1Out_reg_0__0_ ( .D(s1_linMapOut_0__0_), .CK(clk), .Q(
        stage1Out[0]), .QN() );
  DFF_X1 s1_stage1Out_reg_0__1_ ( .D(s1_linMapOut_0__1_), .CK(clk), .Q(
        stage1Out[1]), .QN() );
  DFF_X1 s1_stage1Out_reg_0__2_ ( .D(sboxIn[0]), .CK(clk), .Q(stage1Out[2]), 
        .QN() );
  DFF_X1 s1_stage1Out_reg_0__3_ ( .D(s1_linMapOut_0__3_), .CK(clk), .Q(
        stage1Out[3]), .QN() );
  DFF_X1 s1_stage1Out_reg_0__4_ ( .D(s1_linMapOut_0__4_), .CK(clk), .Q(
        stage1Out[4]), .QN() );
  DFF_X1 s1_stage1Out_reg_0__5_ ( .D(s1_linMapOut_0__5_), .CK(clk), .Q(
        stage1Out[5]), .QN() );
  DFF_X1 s1_stage1Out_reg_0__6_ ( .D(s1_linMapOut_0__6_), .CK(clk), .Q(
        stage1Out[6]), .QN() );
  DFF_X1 s1_stage1Out_reg_0__7_ ( .D(s1_linMapOut_0__7_), .CK(clk), .Q(
        stage1Out[7]), .QN() );
  DFF_X1 s1_stage1Out_reg_1__0_ ( .D(s1_linMapOut_1__0_), .CK(clk), .Q(
        stage1Out[8]), .QN() );
  DFF_X1 s1_stage1Out_reg_1__1_ ( .D(s1_linMapOut_1__1_), .CK(clk), .Q(
        stage1Out[9]), .QN() );
  DFF_X1 s1_stage1Out_reg_1__2_ ( .D(sboxIn[8]), .CK(clk), .Q(stage1Out[10]), 
        .QN() );
  DFF_X1 s1_stage1Out_reg_1__3_ ( .D(s1_linMapOut_1__3_), .CK(clk), .Q(
        stage1Out[11]), .QN() );
  DFF_X1 s1_stage1Out_reg_1__4_ ( .D(s1_linMapOut_1__4_), .CK(clk), .Q(
        stage1Out[12]), .QN() );
  DFF_X1 s1_stage1Out_reg_1__5_ ( .D(s1_linMapOut_1__5_), .CK(clk), .Q(
        stage1Out[13]), .QN() );
  DFF_X1 s1_stage1Out_reg_1__6_ ( .D(s1_linMapOut_1__6_), .CK(clk), .Q(
        stage1Out[14]), .QN() );
  DFF_X1 s1_stage1Out_reg_1__7_ ( .D(s1_linMapOut_1__7_), .CK(clk), .Q(
        stage1Out[15]), .QN() );
  XNOR2_X1 s1_input_mapping_1_U14 ( .A(s1_input_mapping_1_n23), .B(
        s1_input_mapping_1_n22), .ZN(s1_linMapOut_1__7_) );
  XOR2_X1 s1_input_mapping_1_U13 ( .A(sboxIn[12]), .B(s1_linMapOut_1__1_), .Z(
        s1_linMapOut_1__6_) );
  XNOR2_X1 s1_input_mapping_1_U12 ( .A(s1_input_mapping_1_n21), .B(
        s1_input_mapping_1_n20), .ZN(s1_linMapOut_1__5_) );
  XNOR2_X1 s1_input_mapping_1_U11 ( .A(sboxIn[8]), .B(s1_input_mapping_1_n22), 
        .ZN(s1_linMapOut_1__4_) );
  XNOR2_X1 s1_input_mapping_1_U10 ( .A(sboxIn[15]), .B(s1_input_mapping_1_n21), 
        .ZN(s1_input_mapping_1_n22) );
  XNOR2_X1 s1_input_mapping_1_U9 ( .A(s1_input_mapping_1_n19), .B(
        s1_input_mapping_1_n18), .ZN(s1_linMapOut_1__3_) );
  XNOR2_X1 s1_input_mapping_1_U8 ( .A(s1_input_mapping_1_n20), .B(sboxIn[11]), 
        .ZN(s1_input_mapping_1_n18) );
  XNOR2_X1 s1_input_mapping_1_U7 ( .A(sboxIn[15]), .B(sboxIn[12]), .ZN(
        s1_input_mapping_1_n19) );
  XOR2_X1 s1_input_mapping_1_U6 ( .A(sboxIn[8]), .B(s1_input_mapping_1_n21), 
        .Z(s1_linMapOut_1__1_) );
  XOR2_X1 s1_input_mapping_1_U5 ( .A(sboxIn[14]), .B(sboxIn[13]), .Z(
        s1_input_mapping_1_n21) );
  XNOR2_X1 s1_input_mapping_1_U4 ( .A(s1_input_mapping_1_n23), .B(
        s1_input_mapping_1_n17), .ZN(s1_linMapOut_1__0_) );
  XNOR2_X1 s1_input_mapping_1_U3 ( .A(sboxIn[14]), .B(sboxIn[11]), .ZN(
        s1_input_mapping_1_n17) );
  XNOR2_X1 s1_input_mapping_1_U2 ( .A(sboxIn[10]), .B(s1_input_mapping_1_n20), 
        .ZN(s1_input_mapping_1_n23) );
  XNOR2_X1 s1_input_mapping_1_U1 ( .A(sboxIn[8]), .B(sboxIn[9]), .ZN(
        s1_input_mapping_1_n20) );
  XNOR2_X1 s1_input_mapping_0_U14 ( .A(s1_input_mapping_0_n23), .B(
        s1_input_mapping_0_n22), .ZN(s1_linMapOut_0__7_) );
  XOR2_X1 s1_input_mapping_0_U13 ( .A(sboxIn[4]), .B(s1_linMapOut_0__1_), .Z(
        s1_linMapOut_0__6_) );
  XNOR2_X1 s1_input_mapping_0_U12 ( .A(s1_input_mapping_0_n21), .B(
        s1_input_mapping_0_n20), .ZN(s1_linMapOut_0__5_) );
  XNOR2_X1 s1_input_mapping_0_U11 ( .A(sboxIn[0]), .B(s1_input_mapping_0_n22), 
        .ZN(s1_linMapOut_0__4_) );
  XNOR2_X1 s1_input_mapping_0_U10 ( .A(sboxIn[7]), .B(s1_input_mapping_0_n21), 
        .ZN(s1_input_mapping_0_n22) );
  XNOR2_X1 s1_input_mapping_0_U9 ( .A(s1_input_mapping_0_n19), .B(
        s1_input_mapping_0_n18), .ZN(s1_linMapOut_0__3_) );
  XNOR2_X1 s1_input_mapping_0_U8 ( .A(s1_input_mapping_0_n20), .B(sboxIn[3]), 
        .ZN(s1_input_mapping_0_n18) );
  XNOR2_X1 s1_input_mapping_0_U7 ( .A(sboxIn[7]), .B(sboxIn[4]), .ZN(
        s1_input_mapping_0_n19) );
  XOR2_X1 s1_input_mapping_0_U6 ( .A(sboxIn[0]), .B(s1_input_mapping_0_n21), 
        .Z(s1_linMapOut_0__1_) );
  XOR2_X1 s1_input_mapping_0_U5 ( .A(sboxIn[6]), .B(sboxIn[5]), .Z(
        s1_input_mapping_0_n21) );
  XNOR2_X1 s1_input_mapping_0_U4 ( .A(s1_input_mapping_0_n23), .B(
        s1_input_mapping_0_n17), .ZN(s1_linMapOut_0__0_) );
  XNOR2_X1 s1_input_mapping_0_U3 ( .A(sboxIn[6]), .B(sboxIn[3]), .ZN(
        s1_input_mapping_0_n17) );
  XNOR2_X1 s1_input_mapping_0_U2 ( .A(sboxIn[2]), .B(s1_input_mapping_0_n20), 
        .ZN(s1_input_mapping_0_n23) );
  XNOR2_X1 s1_input_mapping_0_U1 ( .A(sboxIn[0]), .B(sboxIn[1]), .ZN(
        s1_input_mapping_0_n20) );
  XOR2_X1 s2_U42 ( .A(stage1Out[11]), .B(stage1Out[15]), .Z(s2_sqsc_in_1__3_)
         );
  XOR2_X1 s2_U41 ( .A(stage1Out[10]), .B(stage1Out[14]), .Z(s2_sqsc_in_1__2_)
         );
  XOR2_X1 s2_U40 ( .A(stage1Out[9]), .B(stage1Out[13]), .Z(s2_sqsc_in_1__1_)
         );
  XOR2_X1 s2_U39 ( .A(stage1Out[3]), .B(stage1Out[7]), .Z(s2_sqsc_in_0__3_) );
  XOR2_X1 s2_U38 ( .A(stage1Out[2]), .B(stage1Out[6]), .Z(s2_sqsc_in_0__2_) );
  XOR2_X1 s2_U37 ( .A(stage1Out[1]), .B(stage1Out[5]), .Z(s2_sqsc_in_0__1_) );
  XOR2_X1 s2_U36 ( .A(s2_sqsc_out[5]), .B(s2_n16), .Z(s2_refreshed[15]) );
  XNOR2_X1 s2_U35 ( .A(s2_n15), .B(s2_n14), .ZN(s2_n16) );
  XNOR2_X1 s2_U34 ( .A(randomS2[7]), .B(randomS2[3]), .ZN(s2_n14) );
  XOR2_X1 s2_U33 ( .A(s2_gf2_mul_out_1__1__3_), .B(randomS2[11]), .Z(s2_n15)
         );
  XOR2_X1 s2_U32 ( .A(s2_sqsc_out[4]), .B(s2_n13), .Z(s2_refreshed[14]) );
  XNOR2_X1 s2_U31 ( .A(s2_n12), .B(s2_n11), .ZN(s2_n13) );
  XNOR2_X1 s2_U30 ( .A(randomS2[6]), .B(randomS2[2]), .ZN(s2_n11) );
  XOR2_X1 s2_U29 ( .A(s2_gf2_mul_out_1__1__2_), .B(randomS2[10]), .Z(s2_n12)
         );
  XOR2_X1 s2_U28 ( .A(s2_sqsc_out[3]), .B(s2_n10), .Z(s2_refreshed[13]) );
  XNOR2_X1 s2_U27 ( .A(s2_n9), .B(s2_n8), .ZN(s2_n10) );
  XNOR2_X1 s2_U26 ( .A(randomS2[5]), .B(randomS2[1]), .ZN(s2_n8) );
  XOR2_X1 s2_U25 ( .A(s2_gf2_mul_out_1__1__1_), .B(randomS2[9]), .Z(s2_n9) );
  XOR2_X1 s2_U24 ( .A(s2_sqsc_in_1__0_), .B(s2_n7), .Z(s2_refreshed[12]) );
  XNOR2_X1 s2_U23 ( .A(s2_n6), .B(s2_n5), .ZN(s2_n7) );
  XNOR2_X1 s2_U22 ( .A(randomS2[8]), .B(randomS2[0]), .ZN(s2_n5) );
  XOR2_X1 s2_U21 ( .A(s2_gf2_mul_out_1__1__0_), .B(randomS2[4]), .Z(s2_n6) );
  XOR2_X1 s2_U20 ( .A(stage1Out[8]), .B(stage1Out[12]), .Z(s2_sqsc_in_1__0_)
         );
  XOR2_X1 s2_U19 ( .A(randomS2[11]), .B(s2_xorResult[7]), .Z(s2_refreshed[11])
         );
  XOR2_X1 s2_U18 ( .A(randomS2[10]), .B(s2_xorResult[6]), .Z(s2_refreshed[10])
         );
  XOR2_X1 s2_U17 ( .A(randomS2[9]), .B(s2_xorResult[5]), .Z(s2_refreshed[9])
         );
  XOR2_X1 s2_U16 ( .A(randomS2[8]), .B(s2_xorResult[4]), .Z(s2_refreshed[8])
         );
  XOR2_X1 s2_U15 ( .A(randomS2[7]), .B(s2_xorResult[3]), .Z(s2_refreshed[7])
         );
  XOR2_X1 s2_U14 ( .A(randomS2[6]), .B(s2_xorResult[2]), .Z(s2_refreshed[6])
         );
  XOR2_X1 s2_U13 ( .A(randomS2[5]), .B(s2_xorResult[1]), .Z(s2_refreshed[5])
         );
  XOR2_X1 s2_U12 ( .A(randomS2[4]), .B(s2_xorResult[0]), .Z(s2_refreshed[4])
         );
  XNOR2_X1 s2_U11 ( .A(s2_n4), .B(s2_sqsc_out[2]), .ZN(s2_refreshed[3]) );
  XNOR2_X1 s2_U10 ( .A(randomS2[3]), .B(s2_gf2_mul_out_0__0__3_), .ZN(s2_n4)
         );
  XNOR2_X1 s2_U9 ( .A(s2_n3), .B(s2_sqsc_out[1]), .ZN(s2_refreshed[2]) );
  XNOR2_X1 s2_U8 ( .A(randomS2[2]), .B(s2_gf2_mul_out_0__0__2_), .ZN(s2_n3) );
  XNOR2_X1 s2_U7 ( .A(s2_n2), .B(s2_sqsc_out[0]), .ZN(s2_refreshed[1]) );
  XNOR2_X1 s2_U6 ( .A(randomS2[1]), .B(s2_gf2_mul_out_0__0__1_), .ZN(s2_n2) );
  XNOR2_X1 s2_U5 ( .A(s2_n1), .B(s2_gf2_mul_out_0__0__0_), .ZN(s2_refreshed[0]) );
  XNOR2_X1 s2_U4 ( .A(randomS2[0]), .B(s2_sqsc_in_0__0_), .ZN(s2_n1) );
  XOR2_X1 s2_U3 ( .A(stage1Out[0]), .B(stage1Out[4]), .Z(s2_sqsc_in_0__0_) );
  DFF_X1 s2_regOut_reg_0__0__0_ ( .D(stage1Out[0]), .CK(clk), .Q(stage2Out[0]), 
        .QN() );
  DFF_X1 s2_regOut_reg_0__0__1_ ( .D(stage1Out[1]), .CK(clk), .Q(stage2Out[1]), 
        .QN() );
  DFF_X1 s2_regOut_reg_0__0__2_ ( .D(stage1Out[2]), .CK(clk), .Q(stage2Out[2]), 
        .QN() );
  DFF_X1 s2_regOut_reg_0__0__3_ ( .D(stage1Out[3]), .CK(clk), .Q(stage2Out[3]), 
        .QN() );
  DFF_X1 s2_regOut_reg_0__1__0_ ( .D(s2_refreshed[0]), .CK(clk), .Q(
        s2_regOut_0__1__0_), .QN() );
  DFF_X1 s2_regOut_reg_0__1__1_ ( .D(s2_refreshed[1]), .CK(clk), .Q(
        s2_regOut_0__1__1_), .QN() );
  DFF_X1 s2_regOut_reg_0__1__2_ ( .D(s2_refreshed[2]), .CK(clk), .Q(
        s2_regOut_0__1__2_), .QN() );
  DFF_X1 s2_regOut_reg_0__1__3_ ( .D(s2_refreshed[3]), .CK(clk), .Q(
        s2_regOut_0__1__3_), .QN() );
  DFF_X1 s2_regOut_reg_0__2__0_ ( .D(s2_refreshed[4]), .CK(clk), .Q(
        s2_regOut_0__2__0_), .QN() );
  DFF_X1 s2_regOut_reg_0__2__1_ ( .D(s2_refreshed[5]), .CK(clk), .Q(
        s2_regOut_0__2__1_), .QN() );
  DFF_X1 s2_regOut_reg_0__2__2_ ( .D(s2_refreshed[6]), .CK(clk), .Q(
        s2_regOut_0__2__2_), .QN() );
  DFF_X1 s2_regOut_reg_0__2__3_ ( .D(s2_refreshed[7]), .CK(clk), .Q(
        s2_regOut_0__2__3_), .QN() );
  DFF_X1 s2_regOut_reg_0__3__0_ ( .D(stage1Out[4]), .CK(clk), .Q(stage2Out[8]), 
        .QN() );
  DFF_X1 s2_regOut_reg_0__3__1_ ( .D(stage1Out[5]), .CK(clk), .Q(stage2Out[9]), 
        .QN() );
  DFF_X1 s2_regOut_reg_0__3__2_ ( .D(stage1Out[6]), .CK(clk), .Q(stage2Out[10]), .QN() );
  DFF_X1 s2_regOut_reg_0__3__3_ ( .D(stage1Out[7]), .CK(clk), .Q(stage2Out[11]), .QN() );
  DFF_X1 s2_regOut_reg_1__0__0_ ( .D(stage1Out[8]), .CK(clk), .Q(stage2Out[12]), .QN() );
  DFF_X1 s2_regOut_reg_1__0__1_ ( .D(stage1Out[9]), .CK(clk), .Q(stage2Out[13]), .QN() );
  DFF_X1 s2_regOut_reg_1__0__2_ ( .D(stage1Out[10]), .CK(clk), .Q(
        stage2Out[14]), .QN() );
  DFF_X1 s2_regOut_reg_1__0__3_ ( .D(stage1Out[11]), .CK(clk), .Q(
        stage2Out[15]), .QN() );
  DFF_X1 s2_regOut_reg_1__1__0_ ( .D(s2_refreshed[8]), .CK(clk), .Q(
        s2_regOut_1__1__0_), .QN() );
  DFF_X1 s2_regOut_reg_1__1__1_ ( .D(s2_refreshed[9]), .CK(clk), .Q(
        s2_regOut_1__1__1_), .QN() );
  DFF_X1 s2_regOut_reg_1__1__2_ ( .D(s2_refreshed[10]), .CK(clk), .Q(
        s2_regOut_1__1__2_), .QN() );
  DFF_X1 s2_regOut_reg_1__1__3_ ( .D(s2_refreshed[11]), .CK(clk), .Q(
        s2_regOut_1__1__3_), .QN() );
  DFF_X1 s2_regOut_reg_1__2__0_ ( .D(s2_refreshed[12]), .CK(clk), .Q(
        s2_regOut_1__2__0_), .QN() );
  DFF_X1 s2_regOut_reg_1__2__1_ ( .D(s2_refreshed[13]), .CK(clk), .Q(
        s2_regOut_1__2__1_), .QN() );
  DFF_X1 s2_regOut_reg_1__2__2_ ( .D(s2_refreshed[14]), .CK(clk), .Q(
        s2_regOut_1__2__2_), .QN() );
  DFF_X1 s2_regOut_reg_1__2__3_ ( .D(s2_refreshed[15]), .CK(clk), .Q(
        s2_regOut_1__2__3_), .QN() );
  DFF_X1 s2_regOut_reg_1__3__0_ ( .D(stage1Out[12]), .CK(clk), .Q(
        stage2Out[20]), .QN() );
  DFF_X1 s2_regOut_reg_1__3__1_ ( .D(stage1Out[13]), .CK(clk), .Q(
        stage2Out[21]), .QN() );
  DFF_X1 s2_regOut_reg_1__3__2_ ( .D(stage1Out[14]), .CK(clk), .Q(
        stage2Out[22]), .QN() );
  DFF_X1 s2_regOut_reg_1__3__3_ ( .D(stage1Out[15]), .CK(clk), .Q(
        stage2Out[23]), .QN() );
  XOR2_X1 s2_sqsc_1_U3 ( .A(s2_sqsc_in_1__0_), .B(s2_sqsc_in_1__2_), .Z(
        s2_sqsc_out[5]) );
  XOR2_X1 s2_sqsc_1_U2 ( .A(s2_sqsc_in_1__1_), .B(s2_sqsc_in_1__3_), .Z(
        s2_sqsc_out[4]) );
  XOR2_X1 s2_sqsc_1_U1 ( .A(s2_sqsc_in_1__0_), .B(s2_sqsc_in_1__1_), .Z(
        s2_sqsc_out[3]) );
  XOR2_X1 s2_sqsc_0_U3 ( .A(s2_sqsc_in_0__0_), .B(s2_sqsc_in_0__2_), .Z(
        s2_sqsc_out[2]) );
  XOR2_X1 s2_sqsc_0_U2 ( .A(s2_sqsc_in_0__1_), .B(s2_sqsc_in_0__3_), .Z(
        s2_sqsc_out[1]) );
  XOR2_X1 s2_sqsc_0_U1 ( .A(s2_sqsc_in_0__0_), .B(s2_sqsc_in_0__1_), .Z(
        s2_sqsc_out[0]) );
  XNOR2_X1 s2_mul1_1_1_U29 ( .A(s2_mul1_1_1_n77), .B(s2_mul1_1_1_n76), .ZN(
        s2_gf2_mul_out_1__1__3_) );
  NAND2_X1 s2_mul1_1_1_U28 ( .A1(stage1Out[15]), .A2(stage1Out[11]), .ZN(
        s2_mul1_1_1_n76) );
  XOR2_X1 s2_mul1_1_1_U27 ( .A(s2_mul1_1_1_n75), .B(s2_mul1_1_1_n74), .Z(
        s2_mul1_1_1_n77) );
  XNOR2_X1 s2_mul1_1_1_U26 ( .A(s2_mul1_1_1_n73), .B(s2_mul1_1_1_n72), .ZN(
        s2_gf2_mul_out_1__1__2_) );
  NAND2_X1 s2_mul1_1_1_U25 ( .A1(stage1Out[14]), .A2(stage1Out[10]), .ZN(
        s2_mul1_1_1_n72) );
  XOR2_X1 s2_mul1_1_1_U24 ( .A(s2_mul1_1_1_n74), .B(s2_mul1_1_1_n71), .Z(
        s2_mul1_1_1_n73) );
  NOR2_X1 s2_mul1_1_1_U23 ( .A1(s2_mul1_1_1_n70), .A2(s2_mul1_1_1_n69), .ZN(
        s2_mul1_1_1_n74) );
  XNOR2_X1 s2_mul1_1_1_U22 ( .A(stage1Out[14]), .B(stage1Out[15]), .ZN(
        s2_mul1_1_1_n69) );
  XNOR2_X1 s2_mul1_1_1_U21 ( .A(stage1Out[10]), .B(stage1Out[11]), .ZN(
        s2_mul1_1_1_n70) );
  XNOR2_X1 s2_mul1_1_1_U20 ( .A(s2_mul1_1_1_n68), .B(s2_mul1_1_1_n67), .ZN(
        s2_gf2_mul_out_1__1__1_) );
  NAND2_X1 s2_mul1_1_1_U19 ( .A1(stage1Out[13]), .A2(stage1Out[9]), .ZN(
        s2_mul1_1_1_n67) );
  XOR2_X1 s2_mul1_1_1_U18 ( .A(s2_mul1_1_1_n75), .B(s2_mul1_1_1_n66), .Z(
        s2_mul1_1_1_n68) );
  XNOR2_X1 s2_mul1_1_1_U17 ( .A(s2_mul1_1_1_n65), .B(s2_mul1_1_1_n64), .ZN(
        s2_mul1_1_1_n75) );
  NAND2_X1 s2_mul1_1_1_U16 ( .A1(s2_mul1_1_1_n63), .A2(s2_mul1_1_1_n62), .ZN(
        s2_mul1_1_1_n64) );
  XNOR2_X1 s2_mul1_1_1_U15 ( .A(s2_mul1_1_1_n61), .B(s2_mul1_1_1_n60), .ZN(
        s2_mul1_1_1_n62) );
  XNOR2_X1 s2_mul1_1_1_U14 ( .A(s2_mul1_1_1_n59), .B(s2_mul1_1_1_n58), .ZN(
        s2_mul1_1_1_n63) );
  XNOR2_X1 s2_mul1_1_1_U13 ( .A(s2_mul1_1_1_n57), .B(s2_mul1_1_1_n56), .ZN(
        s2_gf2_mul_out_1__1__0_) );
  NAND2_X1 s2_mul1_1_1_U12 ( .A1(stage1Out[12]), .A2(stage1Out[8]), .ZN(
        s2_mul1_1_1_n56) );
  XOR2_X1 s2_mul1_1_1_U11 ( .A(s2_mul1_1_1_n66), .B(s2_mul1_1_1_n71), .Z(
        s2_mul1_1_1_n57) );
  XNOR2_X1 s2_mul1_1_1_U10 ( .A(s2_mul1_1_1_n55), .B(s2_mul1_1_1_n65), .ZN(
        s2_mul1_1_1_n71) );
  NOR2_X1 s2_mul1_1_1_U9 ( .A1(s2_mul1_1_1_n61), .A2(s2_mul1_1_1_n59), .ZN(
        s2_mul1_1_1_n65) );
  XNOR2_X1 s2_mul1_1_1_U8 ( .A(stage1Out[12]), .B(stage1Out[14]), .ZN(
        s2_mul1_1_1_n59) );
  XNOR2_X1 s2_mul1_1_1_U7 ( .A(stage1Out[8]), .B(stage1Out[10]), .ZN(
        s2_mul1_1_1_n61) );
  NAND2_X1 s2_mul1_1_1_U6 ( .A1(s2_mul1_1_1_n58), .A2(s2_mul1_1_1_n60), .ZN(
        s2_mul1_1_1_n55) );
  XOR2_X1 s2_mul1_1_1_U5 ( .A(stage1Out[9]), .B(stage1Out[11]), .Z(
        s2_mul1_1_1_n60) );
  XOR2_X1 s2_mul1_1_1_U4 ( .A(stage1Out[13]), .B(stage1Out[15]), .Z(
        s2_mul1_1_1_n58) );
  NOR2_X1 s2_mul1_1_1_U3 ( .A1(s2_mul1_1_1_n54), .A2(s2_mul1_1_1_n53), .ZN(
        s2_mul1_1_1_n66) );
  XNOR2_X1 s2_mul1_1_1_U2 ( .A(stage1Out[12]), .B(stage1Out[13]), .ZN(
        s2_mul1_1_1_n53) );
  XNOR2_X1 s2_mul1_1_1_U1 ( .A(stage1Out[8]), .B(stage1Out[9]), .ZN(
        s2_mul1_1_1_n54) );
  XNOR2_X1 s2_mul1_1_0_U29 ( .A(s2_mul1_1_0_n77), .B(s2_mul1_1_0_n76), .ZN(
        s2_xorResult[7]) );
  NAND2_X1 s2_mul1_1_0_U28 ( .A1(stage1Out[15]), .A2(stage1Out[3]), .ZN(
        s2_mul1_1_0_n76) );
  XOR2_X1 s2_mul1_1_0_U27 ( .A(s2_mul1_1_0_n75), .B(s2_mul1_1_0_n74), .Z(
        s2_mul1_1_0_n77) );
  XNOR2_X1 s2_mul1_1_0_U26 ( .A(s2_mul1_1_0_n73), .B(s2_mul1_1_0_n72), .ZN(
        s2_xorResult[6]) );
  NAND2_X1 s2_mul1_1_0_U25 ( .A1(stage1Out[14]), .A2(stage1Out[2]), .ZN(
        s2_mul1_1_0_n72) );
  XOR2_X1 s2_mul1_1_0_U24 ( .A(s2_mul1_1_0_n74), .B(s2_mul1_1_0_n71), .Z(
        s2_mul1_1_0_n73) );
  NOR2_X1 s2_mul1_1_0_U23 ( .A1(s2_mul1_1_0_n70), .A2(s2_mul1_1_0_n69), .ZN(
        s2_mul1_1_0_n74) );
  XNOR2_X1 s2_mul1_1_0_U22 ( .A(stage1Out[14]), .B(stage1Out[15]), .ZN(
        s2_mul1_1_0_n69) );
  XNOR2_X1 s2_mul1_1_0_U21 ( .A(stage1Out[2]), .B(stage1Out[3]), .ZN(
        s2_mul1_1_0_n70) );
  XNOR2_X1 s2_mul1_1_0_U20 ( .A(s2_mul1_1_0_n68), .B(s2_mul1_1_0_n67), .ZN(
        s2_xorResult[5]) );
  NAND2_X1 s2_mul1_1_0_U19 ( .A1(stage1Out[13]), .A2(stage1Out[1]), .ZN(
        s2_mul1_1_0_n67) );
  XOR2_X1 s2_mul1_1_0_U18 ( .A(s2_mul1_1_0_n75), .B(s2_mul1_1_0_n66), .Z(
        s2_mul1_1_0_n68) );
  XNOR2_X1 s2_mul1_1_0_U17 ( .A(s2_mul1_1_0_n65), .B(s2_mul1_1_0_n64), .ZN(
        s2_mul1_1_0_n75) );
  NAND2_X1 s2_mul1_1_0_U16 ( .A1(s2_mul1_1_0_n63), .A2(s2_mul1_1_0_n62), .ZN(
        s2_mul1_1_0_n64) );
  XNOR2_X1 s2_mul1_1_0_U15 ( .A(s2_mul1_1_0_n61), .B(s2_mul1_1_0_n60), .ZN(
        s2_mul1_1_0_n62) );
  XNOR2_X1 s2_mul1_1_0_U14 ( .A(s2_mul1_1_0_n59), .B(s2_mul1_1_0_n58), .ZN(
        s2_mul1_1_0_n63) );
  XNOR2_X1 s2_mul1_1_0_U13 ( .A(s2_mul1_1_0_n57), .B(s2_mul1_1_0_n56), .ZN(
        s2_xorResult[4]) );
  NAND2_X1 s2_mul1_1_0_U12 ( .A1(stage1Out[12]), .A2(stage1Out[0]), .ZN(
        s2_mul1_1_0_n56) );
  XOR2_X1 s2_mul1_1_0_U11 ( .A(s2_mul1_1_0_n66), .B(s2_mul1_1_0_n71), .Z(
        s2_mul1_1_0_n57) );
  XNOR2_X1 s2_mul1_1_0_U10 ( .A(s2_mul1_1_0_n55), .B(s2_mul1_1_0_n65), .ZN(
        s2_mul1_1_0_n71) );
  NOR2_X1 s2_mul1_1_0_U9 ( .A1(s2_mul1_1_0_n61), .A2(s2_mul1_1_0_n59), .ZN(
        s2_mul1_1_0_n65) );
  XNOR2_X1 s2_mul1_1_0_U8 ( .A(stage1Out[12]), .B(stage1Out[14]), .ZN(
        s2_mul1_1_0_n59) );
  XNOR2_X1 s2_mul1_1_0_U7 ( .A(stage1Out[0]), .B(stage1Out[2]), .ZN(
        s2_mul1_1_0_n61) );
  NAND2_X1 s2_mul1_1_0_U6 ( .A1(s2_mul1_1_0_n58), .A2(s2_mul1_1_0_n60), .ZN(
        s2_mul1_1_0_n55) );
  XOR2_X1 s2_mul1_1_0_U5 ( .A(stage1Out[1]), .B(stage1Out[3]), .Z(
        s2_mul1_1_0_n60) );
  XOR2_X1 s2_mul1_1_0_U4 ( .A(stage1Out[13]), .B(stage1Out[15]), .Z(
        s2_mul1_1_0_n58) );
  NOR2_X1 s2_mul1_1_0_U3 ( .A1(s2_mul1_1_0_n54), .A2(s2_mul1_1_0_n53), .ZN(
        s2_mul1_1_0_n66) );
  XNOR2_X1 s2_mul1_1_0_U2 ( .A(stage1Out[12]), .B(stage1Out[13]), .ZN(
        s2_mul1_1_0_n53) );
  XNOR2_X1 s2_mul1_1_0_U1 ( .A(stage1Out[0]), .B(stage1Out[1]), .ZN(
        s2_mul1_1_0_n54) );
  XNOR2_X1 s2_mul1_0_1_U29 ( .A(s2_mul1_0_1_n77), .B(s2_mul1_0_1_n76), .ZN(
        s2_xorResult[3]) );
  NAND2_X1 s2_mul1_0_1_U28 ( .A1(stage1Out[7]), .A2(stage1Out[11]), .ZN(
        s2_mul1_0_1_n76) );
  XOR2_X1 s2_mul1_0_1_U27 ( .A(s2_mul1_0_1_n75), .B(s2_mul1_0_1_n74), .Z(
        s2_mul1_0_1_n77) );
  XNOR2_X1 s2_mul1_0_1_U26 ( .A(s2_mul1_0_1_n73), .B(s2_mul1_0_1_n72), .ZN(
        s2_xorResult[2]) );
  NAND2_X1 s2_mul1_0_1_U25 ( .A1(stage1Out[6]), .A2(stage1Out[10]), .ZN(
        s2_mul1_0_1_n72) );
  XOR2_X1 s2_mul1_0_1_U24 ( .A(s2_mul1_0_1_n74), .B(s2_mul1_0_1_n71), .Z(
        s2_mul1_0_1_n73) );
  NOR2_X1 s2_mul1_0_1_U23 ( .A1(s2_mul1_0_1_n70), .A2(s2_mul1_0_1_n69), .ZN(
        s2_mul1_0_1_n74) );
  XNOR2_X1 s2_mul1_0_1_U22 ( .A(stage1Out[6]), .B(stage1Out[7]), .ZN(
        s2_mul1_0_1_n69) );
  XNOR2_X1 s2_mul1_0_1_U21 ( .A(stage1Out[10]), .B(stage1Out[11]), .ZN(
        s2_mul1_0_1_n70) );
  XNOR2_X1 s2_mul1_0_1_U20 ( .A(s2_mul1_0_1_n68), .B(s2_mul1_0_1_n67), .ZN(
        s2_xorResult[1]) );
  NAND2_X1 s2_mul1_0_1_U19 ( .A1(stage1Out[5]), .A2(stage1Out[9]), .ZN(
        s2_mul1_0_1_n67) );
  XOR2_X1 s2_mul1_0_1_U18 ( .A(s2_mul1_0_1_n75), .B(s2_mul1_0_1_n66), .Z(
        s2_mul1_0_1_n68) );
  XNOR2_X1 s2_mul1_0_1_U17 ( .A(s2_mul1_0_1_n65), .B(s2_mul1_0_1_n64), .ZN(
        s2_mul1_0_1_n75) );
  NAND2_X1 s2_mul1_0_1_U16 ( .A1(s2_mul1_0_1_n63), .A2(s2_mul1_0_1_n62), .ZN(
        s2_mul1_0_1_n64) );
  XNOR2_X1 s2_mul1_0_1_U15 ( .A(s2_mul1_0_1_n61), .B(s2_mul1_0_1_n60), .ZN(
        s2_mul1_0_1_n62) );
  XNOR2_X1 s2_mul1_0_1_U14 ( .A(s2_mul1_0_1_n59), .B(s2_mul1_0_1_n58), .ZN(
        s2_mul1_0_1_n63) );
  XNOR2_X1 s2_mul1_0_1_U13 ( .A(s2_mul1_0_1_n57), .B(s2_mul1_0_1_n56), .ZN(
        s2_xorResult[0]) );
  NAND2_X1 s2_mul1_0_1_U12 ( .A1(stage1Out[4]), .A2(stage1Out[8]), .ZN(
        s2_mul1_0_1_n56) );
  XOR2_X1 s2_mul1_0_1_U11 ( .A(s2_mul1_0_1_n66), .B(s2_mul1_0_1_n71), .Z(
        s2_mul1_0_1_n57) );
  XNOR2_X1 s2_mul1_0_1_U10 ( .A(s2_mul1_0_1_n55), .B(s2_mul1_0_1_n65), .ZN(
        s2_mul1_0_1_n71) );
  NOR2_X1 s2_mul1_0_1_U9 ( .A1(s2_mul1_0_1_n61), .A2(s2_mul1_0_1_n59), .ZN(
        s2_mul1_0_1_n65) );
  XNOR2_X1 s2_mul1_0_1_U8 ( .A(stage1Out[4]), .B(stage1Out[6]), .ZN(
        s2_mul1_0_1_n59) );
  XNOR2_X1 s2_mul1_0_1_U7 ( .A(stage1Out[8]), .B(stage1Out[10]), .ZN(
        s2_mul1_0_1_n61) );
  NAND2_X1 s2_mul1_0_1_U6 ( .A1(s2_mul1_0_1_n58), .A2(s2_mul1_0_1_n60), .ZN(
        s2_mul1_0_1_n55) );
  XOR2_X1 s2_mul1_0_1_U5 ( .A(stage1Out[9]), .B(stage1Out[11]), .Z(
        s2_mul1_0_1_n60) );
  XOR2_X1 s2_mul1_0_1_U4 ( .A(stage1Out[5]), .B(stage1Out[7]), .Z(
        s2_mul1_0_1_n58) );
  NOR2_X1 s2_mul1_0_1_U3 ( .A1(s2_mul1_0_1_n54), .A2(s2_mul1_0_1_n53), .ZN(
        s2_mul1_0_1_n66) );
  XNOR2_X1 s2_mul1_0_1_U2 ( .A(stage1Out[4]), .B(stage1Out[5]), .ZN(
        s2_mul1_0_1_n53) );
  XNOR2_X1 s2_mul1_0_1_U1 ( .A(stage1Out[8]), .B(stage1Out[9]), .ZN(
        s2_mul1_0_1_n54) );
  XNOR2_X1 s2_mul1_0_0_U29 ( .A(s2_mul1_0_0_n77), .B(s2_mul1_0_0_n76), .ZN(
        s2_gf2_mul_out_0__0__3_) );
  NAND2_X1 s2_mul1_0_0_U28 ( .A1(stage1Out[7]), .A2(stage1Out[3]), .ZN(
        s2_mul1_0_0_n76) );
  XOR2_X1 s2_mul1_0_0_U27 ( .A(s2_mul1_0_0_n75), .B(s2_mul1_0_0_n74), .Z(
        s2_mul1_0_0_n77) );
  XNOR2_X1 s2_mul1_0_0_U26 ( .A(s2_mul1_0_0_n73), .B(s2_mul1_0_0_n72), .ZN(
        s2_gf2_mul_out_0__0__2_) );
  NAND2_X1 s2_mul1_0_0_U25 ( .A1(stage1Out[6]), .A2(stage1Out[2]), .ZN(
        s2_mul1_0_0_n72) );
  XOR2_X1 s2_mul1_0_0_U24 ( .A(s2_mul1_0_0_n74), .B(s2_mul1_0_0_n71), .Z(
        s2_mul1_0_0_n73) );
  NOR2_X1 s2_mul1_0_0_U23 ( .A1(s2_mul1_0_0_n70), .A2(s2_mul1_0_0_n69), .ZN(
        s2_mul1_0_0_n74) );
  XNOR2_X1 s2_mul1_0_0_U22 ( .A(stage1Out[6]), .B(stage1Out[7]), .ZN(
        s2_mul1_0_0_n69) );
  XNOR2_X1 s2_mul1_0_0_U21 ( .A(stage1Out[2]), .B(stage1Out[3]), .ZN(
        s2_mul1_0_0_n70) );
  XNOR2_X1 s2_mul1_0_0_U20 ( .A(s2_mul1_0_0_n68), .B(s2_mul1_0_0_n67), .ZN(
        s2_gf2_mul_out_0__0__1_) );
  NAND2_X1 s2_mul1_0_0_U19 ( .A1(stage1Out[5]), .A2(stage1Out[1]), .ZN(
        s2_mul1_0_0_n67) );
  XOR2_X1 s2_mul1_0_0_U18 ( .A(s2_mul1_0_0_n75), .B(s2_mul1_0_0_n66), .Z(
        s2_mul1_0_0_n68) );
  XNOR2_X1 s2_mul1_0_0_U17 ( .A(s2_mul1_0_0_n65), .B(s2_mul1_0_0_n64), .ZN(
        s2_mul1_0_0_n75) );
  NAND2_X1 s2_mul1_0_0_U16 ( .A1(s2_mul1_0_0_n63), .A2(s2_mul1_0_0_n62), .ZN(
        s2_mul1_0_0_n64) );
  XNOR2_X1 s2_mul1_0_0_U15 ( .A(s2_mul1_0_0_n61), .B(s2_mul1_0_0_n60), .ZN(
        s2_mul1_0_0_n62) );
  XNOR2_X1 s2_mul1_0_0_U14 ( .A(s2_mul1_0_0_n59), .B(s2_mul1_0_0_n58), .ZN(
        s2_mul1_0_0_n63) );
  XNOR2_X1 s2_mul1_0_0_U13 ( .A(s2_mul1_0_0_n57), .B(s2_mul1_0_0_n56), .ZN(
        s2_gf2_mul_out_0__0__0_) );
  NAND2_X1 s2_mul1_0_0_U12 ( .A1(stage1Out[4]), .A2(stage1Out[0]), .ZN(
        s2_mul1_0_0_n56) );
  XOR2_X1 s2_mul1_0_0_U11 ( .A(s2_mul1_0_0_n66), .B(s2_mul1_0_0_n71), .Z(
        s2_mul1_0_0_n57) );
  XNOR2_X1 s2_mul1_0_0_U10 ( .A(s2_mul1_0_0_n55), .B(s2_mul1_0_0_n65), .ZN(
        s2_mul1_0_0_n71) );
  NOR2_X1 s2_mul1_0_0_U9 ( .A1(s2_mul1_0_0_n61), .A2(s2_mul1_0_0_n59), .ZN(
        s2_mul1_0_0_n65) );
  XNOR2_X1 s2_mul1_0_0_U8 ( .A(stage1Out[4]), .B(stage1Out[6]), .ZN(
        s2_mul1_0_0_n59) );
  XNOR2_X1 s2_mul1_0_0_U7 ( .A(stage1Out[0]), .B(stage1Out[2]), .ZN(
        s2_mul1_0_0_n61) );
  NAND2_X1 s2_mul1_0_0_U6 ( .A1(s2_mul1_0_0_n58), .A2(s2_mul1_0_0_n60), .ZN(
        s2_mul1_0_0_n55) );
  XOR2_X1 s2_mul1_0_0_U5 ( .A(stage1Out[1]), .B(stage1Out[3]), .Z(
        s2_mul1_0_0_n60) );
  XOR2_X1 s2_mul1_0_0_U4 ( .A(stage1Out[5]), .B(stage1Out[7]), .Z(
        s2_mul1_0_0_n58) );
  NOR2_X1 s2_mul1_0_0_U3 ( .A1(s2_mul1_0_0_n54), .A2(s2_mul1_0_0_n53), .ZN(
        s2_mul1_0_0_n66) );
  XNOR2_X1 s2_mul1_0_0_U2 ( .A(stage1Out[4]), .B(stage1Out[5]), .ZN(
        s2_mul1_0_0_n53) );
  XNOR2_X1 s2_mul1_0_0_U1 ( .A(stage1Out[0]), .B(stage1Out[1]), .ZN(
        s2_mul1_0_0_n54) );
  XOR2_X1 s2_compr_0_0_U4 ( .A(s2_regOut_0__1__3_), .B(s2_regOut_0__2__3_), 
        .Z(stage2Out[7]) );
  XOR2_X1 s2_compr_0_0_U3 ( .A(s2_regOut_0__1__2_), .B(s2_regOut_0__2__2_), 
        .Z(stage2Out[6]) );
  XOR2_X1 s2_compr_0_0_U2 ( .A(s2_regOut_0__1__1_), .B(s2_regOut_0__2__1_), 
        .Z(stage2Out[5]) );
  XOR2_X1 s2_compr_0_0_U1 ( .A(s2_regOut_0__1__0_), .B(s2_regOut_0__2__0_), 
        .Z(stage2Out[4]) );
  XOR2_X1 s2_compr_1_0_U4 ( .A(s2_regOut_1__1__3_), .B(s2_regOut_1__2__3_), 
        .Z(stage2Out[19]) );
  XOR2_X1 s2_compr_1_0_U3 ( .A(s2_regOut_1__1__2_), .B(s2_regOut_1__2__2_), 
        .Z(stage2Out[18]) );
  XOR2_X1 s2_compr_1_0_U2 ( .A(s2_regOut_1__1__1_), .B(s2_regOut_1__2__1_), 
        .Z(stage2Out[17]) );
  XOR2_X1 s2_compr_1_0_U1 ( .A(s2_regOut_1__1__0_), .B(s2_regOut_1__2__0_), 
        .Z(stage2Out[16]) );
  XOR2_X1 s3_U22 ( .A(stage2Out[16]), .B(stage2Out[18]), .Z(s3_scale_in_1__0_)
         );
  XOR2_X1 s3_U21 ( .A(stage2Out[4]), .B(stage2Out[6]), .Z(s3_scale_in_0__0_)
         );
  XOR2_X1 s3_U20 ( .A(s3_scale_in_1__1_), .B(s3_n8), .Z(s3_refreshed[7]) );
  XNOR2_X1 s3_U19 ( .A(s3_n7), .B(s3_n6), .ZN(s3_n8) );
  XNOR2_X1 s3_U18 ( .A(randomS3[5]), .B(randomS3[1]), .ZN(s3_n6) );
  XOR2_X1 s3_U17 ( .A(s3_gf2_mul_out_1__1__1_), .B(randomS3[3]), .Z(s3_n7) );
  XOR2_X1 s3_U16 ( .A(stage2Out[17]), .B(stage2Out[19]), .Z(s3_scale_in_1__1_)
         );
  XOR2_X1 s3_U15 ( .A(s3_scale_out[1]), .B(s3_n5), .Z(s3_refreshed[6]) );
  XNOR2_X1 s3_U14 ( .A(s3_n4), .B(s3_n3), .ZN(s3_n5) );
  XNOR2_X1 s3_U13 ( .A(randomS3[2]), .B(randomS3[0]), .ZN(s3_n3) );
  XOR2_X1 s3_U12 ( .A(s3_gf2_mul_out_1__1__0_), .B(randomS3[4]), .Z(s3_n4) );
  XOR2_X1 s3_U11 ( .A(randomS3[5]), .B(s3_xorResult[3]), .Z(s3_refreshed[5])
         );
  XOR2_X1 s3_U10 ( .A(randomS3[4]), .B(s3_xorResult[2]), .Z(s3_refreshed[4])
         );
  XOR2_X1 s3_U9 ( .A(randomS3[3]), .B(s3_xorResult[1]), .Z(s3_refreshed[3]) );
  XOR2_X1 s3_U8 ( .A(randomS3[2]), .B(s3_xorResult[0]), .Z(s3_refreshed[2]) );
  XNOR2_X1 s3_U7 ( .A(s3_n2), .B(s3_gf2_mul_out_0__0__1_), .ZN(s3_refreshed[1]) );
  XNOR2_X1 s3_U6 ( .A(randomS3[1]), .B(s3_scale_in_0__1_), .ZN(s3_n2) );
  XOR2_X1 s3_U5 ( .A(stage2Out[5]), .B(stage2Out[7]), .Z(s3_scale_in_0__1_) );
  XNOR2_X1 s3_U4 ( .A(s3_n1), .B(s3_scale_out[0]), .ZN(s3_refreshed[0]) );
  XNOR2_X1 s3_U3 ( .A(randomS3[0]), .B(s3_gf2_mul_out_0__0__0_), .ZN(s3_n1) );
  DFF_X1 s3_regOut_reg_0__0__0_ ( .D(stage2Out[0]), .CK(clk), .Q(stage3Out[0]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__0__1_ ( .D(stage2Out[1]), .CK(clk), .Q(stage3Out[1]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__1__0_ ( .D(stage2Out[2]), .CK(clk), .Q(stage3Out[2]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__1__1_ ( .D(stage2Out[3]), .CK(clk), .Q(stage3Out[3]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__2__0_ ( .D(stage2Out[4]), .CK(clk), .Q(stage3Out[4]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__2__1_ ( .D(stage2Out[5]), .CK(clk), .Q(stage3Out[5]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__3__0_ ( .D(s3_refreshed[0]), .CK(clk), .Q(
        s3_regOut_0__3__0_), .QN() );
  DFF_X1 s3_regOut_reg_0__3__1_ ( .D(s3_refreshed[1]), .CK(clk), .Q(
        s3_regOut_0__3__1_), .QN() );
  DFF_X1 s3_regOut_reg_0__4__0_ ( .D(s3_refreshed[2]), .CK(clk), .Q(
        s3_regOut_0__4__0_), .QN() );
  DFF_X1 s3_regOut_reg_0__4__1_ ( .D(s3_refreshed[3]), .CK(clk), .Q(
        s3_regOut_0__4__1_), .QN() );
  DFF_X1 s3_regOut_reg_0__5__0_ ( .D(stage2Out[6]), .CK(clk), .Q(stage3Out[6]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__5__1_ ( .D(stage2Out[7]), .CK(clk), .Q(stage3Out[7]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__6__0_ ( .D(stage2Out[8]), .CK(clk), .Q(stage3Out[8]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__6__1_ ( .D(stage2Out[9]), .CK(clk), .Q(stage3Out[9]), 
        .QN() );
  DFF_X1 s3_regOut_reg_0__7__0_ ( .D(stage2Out[10]), .CK(clk), .Q(
        stage3Out[10]), .QN() );
  DFF_X1 s3_regOut_reg_0__7__1_ ( .D(stage2Out[11]), .CK(clk), .Q(
        stage3Out[11]), .QN() );
  DFF_X1 s3_regOut_reg_1__0__0_ ( .D(stage2Out[12]), .CK(clk), .Q(
        stage3Out[12]), .QN() );
  DFF_X1 s3_regOut_reg_1__0__1_ ( .D(stage2Out[13]), .CK(clk), .Q(
        stage3Out[13]), .QN() );
  DFF_X1 s3_regOut_reg_1__1__0_ ( .D(stage2Out[14]), .CK(clk), .Q(
        stage3Out[14]), .QN() );
  DFF_X1 s3_regOut_reg_1__1__1_ ( .D(stage2Out[15]), .CK(clk), .Q(
        stage3Out[15]), .QN() );
  DFF_X1 s3_regOut_reg_1__2__0_ ( .D(stage2Out[16]), .CK(clk), .Q(
        stage3Out[16]), .QN() );
  DFF_X1 s3_regOut_reg_1__2__1_ ( .D(stage2Out[17]), .CK(clk), .Q(
        stage3Out[17]), .QN() );
  DFF_X1 s3_regOut_reg_1__3__0_ ( .D(s3_refreshed[4]), .CK(clk), .Q(
        s3_regOut_1__3__0_), .QN() );
  DFF_X1 s3_regOut_reg_1__3__1_ ( .D(s3_refreshed[5]), .CK(clk), .Q(
        s3_regOut_1__3__1_), .QN() );
  DFF_X1 s3_regOut_reg_1__4__0_ ( .D(s3_refreshed[6]), .CK(clk), .Q(
        s3_regOut_1__4__0_), .QN() );
  DFF_X1 s3_regOut_reg_1__4__1_ ( .D(s3_refreshed[7]), .CK(clk), .Q(
        s3_regOut_1__4__1_), .QN() );
  DFF_X1 s3_regOut_reg_1__5__0_ ( .D(stage2Out[18]), .CK(clk), .Q(
        stage3Out[18]), .QN() );
  DFF_X1 s3_regOut_reg_1__5__1_ ( .D(stage2Out[19]), .CK(clk), .Q(
        stage3Out[19]), .QN() );
  DFF_X1 s3_regOut_reg_1__6__0_ ( .D(stage2Out[20]), .CK(clk), .Q(
        stage3Out[20]), .QN() );
  DFF_X1 s3_regOut_reg_1__6__1_ ( .D(stage2Out[21]), .CK(clk), .Q(
        stage3Out[21]), .QN() );
  DFF_X1 s3_regOut_reg_1__7__0_ ( .D(stage2Out[22]), .CK(clk), .Q(
        stage3Out[22]), .QN() );
  DFF_X1 s3_regOut_reg_1__7__1_ ( .D(stage2Out[23]), .CK(clk), .Q(
        stage3Out[23]), .QN() );
  XOR2_X1 s3_sqsc_1_U1 ( .A(s3_scale_in_1__0_), .B(s3_scale_in_1__1_), .Z(
        s3_scale_out[1]) );
  XOR2_X1 s3_sqsc_0_U1 ( .A(s3_scale_in_0__0_), .B(s3_scale_in_0__1_), .Z(
        s3_scale_out[0]) );
  XNOR2_X1 s3_mul1_1_1_U7 ( .A(s3_mul1_1_1_n15), .B(s3_mul1_1_1_n14), .ZN(
        s3_gf2_mul_out_1__1__1_) );
  NAND2_X1 s3_mul1_1_1_U6 ( .A1(stage2Out[19]), .A2(stage2Out[17]), .ZN(
        s3_mul1_1_1_n15) );
  XNOR2_X1 s3_mul1_1_1_U5 ( .A(s3_mul1_1_1_n13), .B(s3_mul1_1_1_n14), .ZN(
        s3_gf2_mul_out_1__1__0_) );
  NOR2_X1 s3_mul1_1_1_U4 ( .A1(s3_mul1_1_1_n12), .A2(s3_mul1_1_1_n11), .ZN(
        s3_mul1_1_1_n14) );
  XNOR2_X1 s3_mul1_1_1_U3 ( .A(stage2Out[19]), .B(stage2Out[18]), .ZN(
        s3_mul1_1_1_n11) );
  XNOR2_X1 s3_mul1_1_1_U2 ( .A(stage2Out[17]), .B(stage2Out[16]), .ZN(
        s3_mul1_1_1_n12) );
  NAND2_X1 s3_mul1_1_1_U1 ( .A1(stage2Out[18]), .A2(stage2Out[16]), .ZN(
        s3_mul1_1_1_n13) );
  XNOR2_X1 s3_mul1_1_0_U7 ( .A(s3_mul1_1_0_n15), .B(s3_mul1_1_0_n14), .ZN(
        s3_xorResult[3]) );
  NAND2_X1 s3_mul1_1_0_U6 ( .A1(stage2Out[19]), .A2(stage2Out[5]), .ZN(
        s3_mul1_1_0_n15) );
  XNOR2_X1 s3_mul1_1_0_U5 ( .A(s3_mul1_1_0_n13), .B(s3_mul1_1_0_n14), .ZN(
        s3_xorResult[2]) );
  NOR2_X1 s3_mul1_1_0_U4 ( .A1(s3_mul1_1_0_n12), .A2(s3_mul1_1_0_n11), .ZN(
        s3_mul1_1_0_n14) );
  XNOR2_X1 s3_mul1_1_0_U3 ( .A(stage2Out[19]), .B(stage2Out[18]), .ZN(
        s3_mul1_1_0_n11) );
  XNOR2_X1 s3_mul1_1_0_U2 ( .A(stage2Out[5]), .B(stage2Out[4]), .ZN(
        s3_mul1_1_0_n12) );
  NAND2_X1 s3_mul1_1_0_U1 ( .A1(stage2Out[18]), .A2(stage2Out[4]), .ZN(
        s3_mul1_1_0_n13) );
  XNOR2_X1 s3_mul1_0_1_U7 ( .A(s3_mul1_0_1_n15), .B(s3_mul1_0_1_n14), .ZN(
        s3_xorResult[1]) );
  NAND2_X1 s3_mul1_0_1_U6 ( .A1(stage2Out[7]), .A2(stage2Out[17]), .ZN(
        s3_mul1_0_1_n15) );
  XNOR2_X1 s3_mul1_0_1_U5 ( .A(s3_mul1_0_1_n13), .B(s3_mul1_0_1_n14), .ZN(
        s3_xorResult[0]) );
  NOR2_X1 s3_mul1_0_1_U4 ( .A1(s3_mul1_0_1_n12), .A2(s3_mul1_0_1_n11), .ZN(
        s3_mul1_0_1_n14) );
  XNOR2_X1 s3_mul1_0_1_U3 ( .A(stage2Out[7]), .B(stage2Out[6]), .ZN(
        s3_mul1_0_1_n11) );
  XNOR2_X1 s3_mul1_0_1_U2 ( .A(stage2Out[17]), .B(stage2Out[16]), .ZN(
        s3_mul1_0_1_n12) );
  NAND2_X1 s3_mul1_0_1_U1 ( .A1(stage2Out[6]), .A2(stage2Out[16]), .ZN(
        s3_mul1_0_1_n13) );
  XNOR2_X1 s3_mul1_0_0_U7 ( .A(s3_mul1_0_0_n15), .B(s3_mul1_0_0_n14), .ZN(
        s3_gf2_mul_out_0__0__1_) );
  NAND2_X1 s3_mul1_0_0_U6 ( .A1(stage2Out[7]), .A2(stage2Out[5]), .ZN(
        s3_mul1_0_0_n15) );
  XNOR2_X1 s3_mul1_0_0_U5 ( .A(s3_mul1_0_0_n13), .B(s3_mul1_0_0_n14), .ZN(
        s3_gf2_mul_out_0__0__0_) );
  NOR2_X1 s3_mul1_0_0_U4 ( .A1(s3_mul1_0_0_n12), .A2(s3_mul1_0_0_n11), .ZN(
        s3_mul1_0_0_n14) );
  XNOR2_X1 s3_mul1_0_0_U3 ( .A(stage2Out[7]), .B(stage2Out[6]), .ZN(
        s3_mul1_0_0_n11) );
  XNOR2_X1 s3_mul1_0_0_U2 ( .A(stage2Out[5]), .B(stage2Out[4]), .ZN(
        s3_mul1_0_0_n12) );
  NAND2_X1 s3_mul1_0_0_U1 ( .A1(stage2Out[6]), .A2(stage2Out[4]), .ZN(
        s3_mul1_0_0_n13) );
  XOR2_X1 s3_compr_0_0_U2 ( .A(s3_regOut_0__3__1_), .B(s3_regOut_0__4__1_), 
        .Z(s4_inv_out_0__0_) );
  XOR2_X1 s3_compr_0_0_U1 ( .A(s3_regOut_0__3__0_), .B(s3_regOut_0__4__0_), 
        .Z(s4_inv_out_0__1_) );
  XOR2_X1 s3_compr_1_0_U2 ( .A(s3_regOut_1__3__1_), .B(s3_regOut_1__4__1_), 
        .Z(s4_inv_out_1__0_) );
  XOR2_X1 s3_compr_1_0_U1 ( .A(s3_regOut_1__3__0_), .B(s3_regOut_1__4__0_), 
        .Z(s4_inv_out_1__1_) );
  XNOR2_X1 s4_U26 ( .A(s4_n8), .B(s4_n7), .ZN(s4_refreshed[15]) );
  XNOR2_X1 s4_U25 ( .A(s4_concat[15]), .B(randomS4[11]), .ZN(s4_n7) );
  XOR2_X1 s4_U24 ( .A(randomS4[3]), .B(randomS4[7]), .Z(s4_n8) );
  XNOR2_X1 s4_U23 ( .A(s4_n6), .B(s4_n5), .ZN(s4_refreshed[14]) );
  XNOR2_X1 s4_U22 ( .A(s4_concat[14]), .B(randomS4[10]), .ZN(s4_n5) );
  XOR2_X1 s4_U21 ( .A(randomS4[2]), .B(randomS4[6]), .Z(s4_n6) );
  XNOR2_X1 s4_U20 ( .A(s4_n4), .B(s4_n3), .ZN(s4_refreshed[13]) );
  XNOR2_X1 s4_U19 ( .A(s4_concat[13]), .B(randomS4[9]), .ZN(s4_n3) );
  XOR2_X1 s4_U18 ( .A(randomS4[1]), .B(randomS4[5]), .Z(s4_n4) );
  XNOR2_X1 s4_U17 ( .A(s4_n2), .B(s4_n1), .ZN(s4_refreshed[12]) );
  XNOR2_X1 s4_U16 ( .A(s4_concat[12]), .B(randomS4[8]), .ZN(s4_n1) );
  XOR2_X1 s4_U15 ( .A(randomS4[0]), .B(randomS4[4]), .Z(s4_n2) );
  XOR2_X1 s4_U14 ( .A(randomS4[11]), .B(s4_concat[11]), .Z(s4_refreshed[11])
         );
  XOR2_X1 s4_U13 ( .A(randomS4[10]), .B(s4_concat[10]), .Z(s4_refreshed[10])
         );
  XOR2_X1 s4_U12 ( .A(randomS4[9]), .B(s4_concat[9]), .Z(s4_refreshed[9]) );
  XOR2_X1 s4_U11 ( .A(randomS4[8]), .B(s4_concat[8]), .Z(s4_refreshed[8]) );
  XOR2_X1 s4_U10 ( .A(randomS4[7]), .B(s4_concat[7]), .Z(s4_refreshed[7]) );
  XOR2_X1 s4_U9 ( .A(randomS4[6]), .B(s4_concat[6]), .Z(s4_refreshed[6]) );
  XOR2_X1 s4_U8 ( .A(randomS4[5]), .B(s4_concat[5]), .Z(s4_refreshed[5]) );
  XOR2_X1 s4_U7 ( .A(randomS4[4]), .B(s4_concat[4]), .Z(s4_refreshed[4]) );
  XOR2_X1 s4_U6 ( .A(randomS4[3]), .B(s4_concat[3]), .Z(s4_refreshed[3]) );
  XOR2_X1 s4_U5 ( .A(randomS4[2]), .B(s4_concat[2]), .Z(s4_refreshed[2]) );
  XOR2_X1 s4_U4 ( .A(randomS4[1]), .B(s4_concat[1]), .Z(s4_refreshed[1]) );
  XOR2_X1 s4_U3 ( .A(randomS4[0]), .B(s4_concat[0]), .Z(s4_refreshed[0]) );
  DFF_X1 s4_regOut_reg_0__0__0_ ( .D(stage3Out[0]), .CK(clk), .Q(stage4Out[0]), 
        .QN() );
  DFF_X1 s4_regOut_reg_0__0__1_ ( .D(stage3Out[1]), .CK(clk), .Q(stage4Out[1]), 
        .QN() );
  DFF_X1 s4_regOut_reg_0__0__2_ ( .D(stage3Out[2]), .CK(clk), .Q(stage4Out[2]), 
        .QN() );
  DFF_X1 s4_regOut_reg_0__0__3_ ( .D(stage3Out[3]), .CK(clk), .Q(stage4Out[3]), 
        .QN() );
  DFF_X1 s4_regOut_reg_0__1__0_ ( .D(s4_refreshed[0]), .CK(clk), .Q(
        s4_regOut_0__1__0_), .QN() );
  DFF_X1 s4_regOut_reg_0__1__1_ ( .D(s4_refreshed[1]), .CK(clk), .Q(
        s4_regOut_0__1__1_), .QN() );
  DFF_X1 s4_regOut_reg_0__1__2_ ( .D(s4_refreshed[2]), .CK(clk), .Q(
        s4_regOut_0__1__2_), .QN() );
  DFF_X1 s4_regOut_reg_0__1__3_ ( .D(s4_refreshed[3]), .CK(clk), .Q(
        s4_regOut_0__1__3_), .QN() );
  DFF_X1 s4_regOut_reg_0__2__0_ ( .D(s4_refreshed[4]), .CK(clk), .Q(
        s4_regOut_0__2__0_), .QN() );
  DFF_X1 s4_regOut_reg_0__2__1_ ( .D(s4_refreshed[5]), .CK(clk), .Q(
        s4_regOut_0__2__1_), .QN() );
  DFF_X1 s4_regOut_reg_0__2__2_ ( .D(s4_refreshed[6]), .CK(clk), .Q(
        s4_regOut_0__2__2_), .QN() );
  DFF_X1 s4_regOut_reg_0__2__3_ ( .D(s4_refreshed[7]), .CK(clk), .Q(
        s4_regOut_0__2__3_), .QN() );
  DFF_X1 s4_regOut_reg_0__3__0_ ( .D(stage3Out[8]), .CK(clk), .Q(stage4Out[8]), 
        .QN() );
  DFF_X1 s4_regOut_reg_0__3__1_ ( .D(stage3Out[9]), .CK(clk), .Q(stage4Out[9]), 
        .QN() );
  DFF_X1 s4_regOut_reg_0__3__2_ ( .D(stage3Out[10]), .CK(clk), .Q(
        stage4Out[10]), .QN() );
  DFF_X1 s4_regOut_reg_0__3__3_ ( .D(stage3Out[11]), .CK(clk), .Q(
        stage4Out[11]), .QN() );
  DFF_X1 s4_regOut_reg_1__0__0_ ( .D(stage3Out[12]), .CK(clk), .Q(
        stage4Out[12]), .QN() );
  DFF_X1 s4_regOut_reg_1__0__1_ ( .D(stage3Out[13]), .CK(clk), .Q(
        stage4Out[13]), .QN() );
  DFF_X1 s4_regOut_reg_1__0__2_ ( .D(stage3Out[14]), .CK(clk), .Q(
        stage4Out[14]), .QN() );
  DFF_X1 s4_regOut_reg_1__0__3_ ( .D(stage3Out[15]), .CK(clk), .Q(
        stage4Out[15]), .QN() );
  DFF_X1 s4_regOut_reg_1__1__0_ ( .D(s4_refreshed[8]), .CK(clk), .Q(
        s4_regOut_1__1__0_), .QN() );
  DFF_X1 s4_regOut_reg_1__1__1_ ( .D(s4_refreshed[9]), .CK(clk), .Q(
        s4_regOut_1__1__1_), .QN() );
  DFF_X1 s4_regOut_reg_1__1__2_ ( .D(s4_refreshed[10]), .CK(clk), .Q(
        s4_regOut_1__1__2_), .QN() );
  DFF_X1 s4_regOut_reg_1__1__3_ ( .D(s4_refreshed[11]), .CK(clk), .Q(
        s4_regOut_1__1__3_), .QN() );
  DFF_X1 s4_regOut_reg_1__2__0_ ( .D(s4_refreshed[12]), .CK(clk), .Q(
        s4_regOut_1__2__0_), .QN() );
  DFF_X1 s4_regOut_reg_1__2__1_ ( .D(s4_refreshed[13]), .CK(clk), .Q(
        s4_regOut_1__2__1_), .QN() );
  DFF_X1 s4_regOut_reg_1__2__2_ ( .D(s4_refreshed[14]), .CK(clk), .Q(
        s4_regOut_1__2__2_), .QN() );
  DFF_X1 s4_regOut_reg_1__2__3_ ( .D(s4_refreshed[15]), .CK(clk), .Q(
        s4_regOut_1__2__3_), .QN() );
  DFF_X1 s4_regOut_reg_1__3__0_ ( .D(stage3Out[20]), .CK(clk), .Q(
        stage4Out[20]), .QN() );
  DFF_X1 s4_regOut_reg_1__3__1_ ( .D(stage3Out[21]), .CK(clk), .Q(
        stage4Out[21]), .QN() );
  DFF_X1 s4_regOut_reg_1__3__2_ ( .D(stage3Out[22]), .CK(clk), .Q(
        stage4Out[22]), .QN() );
  DFF_X1 s4_regOut_reg_1__3__3_ ( .D(stage3Out[23]), .CK(clk), .Q(
        stage4Out[23]), .QN() );
  XNOR2_X1 s4_mul1_1_1_U7 ( .A(s4_mul1_1_1_n15), .B(s4_mul1_1_1_n14), .ZN(
        s4_concat[13]) );
  NAND2_X1 s4_mul1_1_1_U6 ( .A1(stage3Out[19]), .A2(s4_inv_out_1__1_), .ZN(
        s4_mul1_1_1_n15) );
  XNOR2_X1 s4_mul1_1_1_U5 ( .A(s4_mul1_1_1_n13), .B(s4_mul1_1_1_n14), .ZN(
        s4_concat[12]) );
  NOR2_X1 s4_mul1_1_1_U4 ( .A1(s4_mul1_1_1_n12), .A2(s4_mul1_1_1_n11), .ZN(
        s4_mul1_1_1_n14) );
  XNOR2_X1 s4_mul1_1_1_U3 ( .A(stage3Out[19]), .B(stage3Out[18]), .ZN(
        s4_mul1_1_1_n11) );
  XNOR2_X1 s4_mul1_1_1_U2 ( .A(s4_inv_out_1__1_), .B(s4_inv_out_1__0_), .ZN(
        s4_mul1_1_1_n12) );
  NAND2_X1 s4_mul1_1_1_U1 ( .A1(stage3Out[18]), .A2(s4_inv_out_1__0_), .ZN(
        s4_mul1_1_1_n13) );
  XNOR2_X1 s4_mul1_1_0_U7 ( .A(s4_mul1_1_0_n15), .B(s4_mul1_1_0_n14), .ZN(
        s4_concat[9]) );
  NAND2_X1 s4_mul1_1_0_U6 ( .A1(stage3Out[19]), .A2(s4_inv_out_0__1_), .ZN(
        s4_mul1_1_0_n15) );
  XNOR2_X1 s4_mul1_1_0_U5 ( .A(s4_mul1_1_0_n13), .B(s4_mul1_1_0_n14), .ZN(
        s4_concat[8]) );
  NOR2_X1 s4_mul1_1_0_U4 ( .A1(s4_mul1_1_0_n12), .A2(s4_mul1_1_0_n11), .ZN(
        s4_mul1_1_0_n14) );
  XNOR2_X1 s4_mul1_1_0_U3 ( .A(stage3Out[19]), .B(stage3Out[18]), .ZN(
        s4_mul1_1_0_n11) );
  XNOR2_X1 s4_mul1_1_0_U2 ( .A(s4_inv_out_0__1_), .B(s4_inv_out_0__0_), .ZN(
        s4_mul1_1_0_n12) );
  NAND2_X1 s4_mul1_1_0_U1 ( .A1(stage3Out[18]), .A2(s4_inv_out_0__0_), .ZN(
        s4_mul1_1_0_n13) );
  XNOR2_X1 s4_mul1_0_1_U7 ( .A(s4_mul1_0_1_n15), .B(s4_mul1_0_1_n14), .ZN(
        s4_concat[5]) );
  NAND2_X1 s4_mul1_0_1_U6 ( .A1(stage3Out[7]), .A2(s4_inv_out_1__1_), .ZN(
        s4_mul1_0_1_n15) );
  XNOR2_X1 s4_mul1_0_1_U5 ( .A(s4_mul1_0_1_n13), .B(s4_mul1_0_1_n14), .ZN(
        s4_concat[4]) );
  NOR2_X1 s4_mul1_0_1_U4 ( .A1(s4_mul1_0_1_n12), .A2(s4_mul1_0_1_n11), .ZN(
        s4_mul1_0_1_n14) );
  XNOR2_X1 s4_mul1_0_1_U3 ( .A(stage3Out[7]), .B(stage3Out[6]), .ZN(
        s4_mul1_0_1_n11) );
  XNOR2_X1 s4_mul1_0_1_U2 ( .A(s4_inv_out_1__1_), .B(s4_inv_out_1__0_), .ZN(
        s4_mul1_0_1_n12) );
  NAND2_X1 s4_mul1_0_1_U1 ( .A1(stage3Out[6]), .A2(s4_inv_out_1__0_), .ZN(
        s4_mul1_0_1_n13) );
  XNOR2_X1 s4_mul1_0_0_U7 ( .A(s4_mul1_0_0_n15), .B(s4_mul1_0_0_n14), .ZN(
        s4_concat[1]) );
  NAND2_X1 s4_mul1_0_0_U6 ( .A1(stage3Out[7]), .A2(s4_inv_out_0__1_), .ZN(
        s4_mul1_0_0_n15) );
  XNOR2_X1 s4_mul1_0_0_U5 ( .A(s4_mul1_0_0_n13), .B(s4_mul1_0_0_n14), .ZN(
        s4_concat[0]) );
  NOR2_X1 s4_mul1_0_0_U4 ( .A1(s4_mul1_0_0_n12), .A2(s4_mul1_0_0_n11), .ZN(
        s4_mul1_0_0_n14) );
  XNOR2_X1 s4_mul1_0_0_U3 ( .A(stage3Out[7]), .B(stage3Out[6]), .ZN(
        s4_mul1_0_0_n11) );
  XNOR2_X1 s4_mul1_0_0_U2 ( .A(s4_inv_out_0__1_), .B(s4_inv_out_0__0_), .ZN(
        s4_mul1_0_0_n12) );
  NAND2_X1 s4_mul1_0_0_U1 ( .A1(stage3Out[6]), .A2(s4_inv_out_0__0_), .ZN(
        s4_mul1_0_0_n13) );
  XNOR2_X1 s4_mul2_1_1_U7 ( .A(s4_mul2_1_1_n15), .B(s4_mul2_1_1_n14), .ZN(
        s4_concat[15]) );
  NAND2_X1 s4_mul2_1_1_U6 ( .A1(stage3Out[17]), .A2(s4_inv_out_1__1_), .ZN(
        s4_mul2_1_1_n15) );
  XNOR2_X1 s4_mul2_1_1_U5 ( .A(s4_mul2_1_1_n13), .B(s4_mul2_1_1_n14), .ZN(
        s4_concat[14]) );
  NOR2_X1 s4_mul2_1_1_U4 ( .A1(s4_mul2_1_1_n12), .A2(s4_mul2_1_1_n11), .ZN(
        s4_mul2_1_1_n14) );
  XNOR2_X1 s4_mul2_1_1_U3 ( .A(stage3Out[17]), .B(stage3Out[16]), .ZN(
        s4_mul2_1_1_n11) );
  XNOR2_X1 s4_mul2_1_1_U2 ( .A(s4_inv_out_1__1_), .B(s4_inv_out_1__0_), .ZN(
        s4_mul2_1_1_n12) );
  NAND2_X1 s4_mul2_1_1_U1 ( .A1(stage3Out[16]), .A2(s4_inv_out_1__0_), .ZN(
        s4_mul2_1_1_n13) );
  XNOR2_X1 s4_mul2_1_0_U7 ( .A(s4_mul2_1_0_n15), .B(s4_mul2_1_0_n14), .ZN(
        s4_concat[11]) );
  NAND2_X1 s4_mul2_1_0_U6 ( .A1(stage3Out[17]), .A2(s4_inv_out_0__1_), .ZN(
        s4_mul2_1_0_n15) );
  XNOR2_X1 s4_mul2_1_0_U5 ( .A(s4_mul2_1_0_n13), .B(s4_mul2_1_0_n14), .ZN(
        s4_concat[10]) );
  NOR2_X1 s4_mul2_1_0_U4 ( .A1(s4_mul2_1_0_n12), .A2(s4_mul2_1_0_n11), .ZN(
        s4_mul2_1_0_n14) );
  XNOR2_X1 s4_mul2_1_0_U3 ( .A(stage3Out[17]), .B(stage3Out[16]), .ZN(
        s4_mul2_1_0_n11) );
  XNOR2_X1 s4_mul2_1_0_U2 ( .A(s4_inv_out_0__1_), .B(s4_inv_out_0__0_), .ZN(
        s4_mul2_1_0_n12) );
  NAND2_X1 s4_mul2_1_0_U1 ( .A1(stage3Out[16]), .A2(s4_inv_out_0__0_), .ZN(
        s4_mul2_1_0_n13) );
  XNOR2_X1 s4_mul2_0_1_U7 ( .A(s4_mul2_0_1_n15), .B(s4_mul2_0_1_n14), .ZN(
        s4_concat[7]) );
  NAND2_X1 s4_mul2_0_1_U6 ( .A1(stage3Out[5]), .A2(s4_inv_out_1__1_), .ZN(
        s4_mul2_0_1_n15) );
  XNOR2_X1 s4_mul2_0_1_U5 ( .A(s4_mul2_0_1_n13), .B(s4_mul2_0_1_n14), .ZN(
        s4_concat[6]) );
  NOR2_X1 s4_mul2_0_1_U4 ( .A1(s4_mul2_0_1_n12), .A2(s4_mul2_0_1_n11), .ZN(
        s4_mul2_0_1_n14) );
  XNOR2_X1 s4_mul2_0_1_U3 ( .A(stage3Out[5]), .B(stage3Out[4]), .ZN(
        s4_mul2_0_1_n11) );
  XNOR2_X1 s4_mul2_0_1_U2 ( .A(s4_inv_out_1__1_), .B(s4_inv_out_1__0_), .ZN(
        s4_mul2_0_1_n12) );
  NAND2_X1 s4_mul2_0_1_U1 ( .A1(stage3Out[4]), .A2(s4_inv_out_1__0_), .ZN(
        s4_mul2_0_1_n13) );
  XNOR2_X1 s4_mul2_0_0_U7 ( .A(s4_mul2_0_0_n15), .B(s4_mul2_0_0_n14), .ZN(
        s4_concat[3]) );
  NAND2_X1 s4_mul2_0_0_U6 ( .A1(stage3Out[5]), .A2(s4_inv_out_0__1_), .ZN(
        s4_mul2_0_0_n15) );
  XNOR2_X1 s4_mul2_0_0_U5 ( .A(s4_mul2_0_0_n13), .B(s4_mul2_0_0_n14), .ZN(
        s4_concat[2]) );
  NOR2_X1 s4_mul2_0_0_U4 ( .A1(s4_mul2_0_0_n12), .A2(s4_mul2_0_0_n11), .ZN(
        s4_mul2_0_0_n14) );
  XNOR2_X1 s4_mul2_0_0_U3 ( .A(stage3Out[5]), .B(stage3Out[4]), .ZN(
        s4_mul2_0_0_n11) );
  XNOR2_X1 s4_mul2_0_0_U2 ( .A(s4_inv_out_0__1_), .B(s4_inv_out_0__0_), .ZN(
        s4_mul2_0_0_n12) );
  NAND2_X1 s4_mul2_0_0_U1 ( .A1(stage3Out[4]), .A2(s4_inv_out_0__0_), .ZN(
        s4_mul2_0_0_n13) );
  XOR2_X2 s4_compr_0_0_U4 ( .A(s4_regOut_0__1__3_), .B(s4_regOut_0__2__3_), 
        .Z(stage4Out[7]) );
  XOR2_X2 s4_compr_0_0_U3 ( .A(s4_regOut_0__1__0_), .B(s4_regOut_0__2__0_), 
        .Z(stage4Out[4]) );
  XOR2_X2 s4_compr_0_0_U2 ( .A(s4_regOut_0__1__2_), .B(s4_regOut_0__2__2_), 
        .Z(stage4Out[6]) );
  XOR2_X2 s4_compr_0_0_U1 ( .A(s4_regOut_0__1__1_), .B(s4_regOut_0__2__1_), 
        .Z(stage4Out[5]) );
  XOR2_X2 s4_compr_1_0_U4 ( .A(s4_regOut_1__1__3_), .B(s4_regOut_1__2__3_), 
        .Z(stage4Out[19]) );
  XOR2_X2 s4_compr_1_0_U3 ( .A(s4_regOut_1__1__0_), .B(s4_regOut_1__2__0_), 
        .Z(stage4Out[16]) );
  XOR2_X2 s4_compr_1_0_U2 ( .A(s4_regOut_1__1__2_), .B(s4_regOut_1__2__2_), 
        .Z(stage4Out[18]) );
  XOR2_X2 s4_compr_1_0_U1 ( .A(s4_regOut_1__1__1_), .B(s4_regOut_1__2__1_), 
        .Z(stage4Out[17]) );
  XNOR2_X1 s5_U50 ( .A(s5_n16), .B(s5_n15), .ZN(s5_refreshed[31]) );
  XNOR2_X1 s5_U49 ( .A(s5_concat[31]), .B(randomS5[23]), .ZN(s5_n15) );
  XOR2_X1 s5_U48 ( .A(randomS5[7]), .B(randomS5[15]), .Z(s5_n16) );
  XNOR2_X1 s5_U47 ( .A(s5_n14), .B(s5_n13), .ZN(s5_refreshed[30]) );
  XNOR2_X1 s5_U46 ( .A(s5_concat[30]), .B(randomS5[22]), .ZN(s5_n13) );
  XOR2_X1 s5_U45 ( .A(randomS5[6]), .B(randomS5[14]), .Z(s5_n14) );
  XNOR2_X1 s5_U44 ( .A(s5_n12), .B(s5_n11), .ZN(s5_refreshed[29]) );
  XNOR2_X1 s5_U43 ( .A(s5_concat[29]), .B(randomS5[21]), .ZN(s5_n11) );
  XOR2_X1 s5_U42 ( .A(randomS5[5]), .B(randomS5[13]), .Z(s5_n12) );
  XNOR2_X1 s5_U41 ( .A(s5_n10), .B(s5_n9), .ZN(s5_refreshed[28]) );
  XNOR2_X1 s5_U40 ( .A(s5_concat[28]), .B(randomS5[20]), .ZN(s5_n9) );
  XOR2_X1 s5_U39 ( .A(randomS5[4]), .B(randomS5[12]), .Z(s5_n10) );
  XNOR2_X1 s5_U38 ( .A(s5_n8), .B(s5_n7), .ZN(s5_refreshed[27]) );
  XNOR2_X1 s5_U37 ( .A(s5_concat[27]), .B(randomS5[19]), .ZN(s5_n7) );
  XOR2_X1 s5_U36 ( .A(randomS5[3]), .B(randomS5[11]), .Z(s5_n8) );
  XNOR2_X1 s5_U35 ( .A(s5_n6), .B(s5_n5), .ZN(s5_refreshed[26]) );
  XNOR2_X1 s5_U34 ( .A(s5_concat[26]), .B(randomS5[18]), .ZN(s5_n5) );
  XOR2_X1 s5_U33 ( .A(randomS5[2]), .B(randomS5[10]), .Z(s5_n6) );
  XNOR2_X1 s5_U32 ( .A(s5_n4), .B(s5_n3), .ZN(s5_refreshed[25]) );
  XNOR2_X1 s5_U31 ( .A(s5_concat[25]), .B(randomS5[17]), .ZN(s5_n3) );
  XOR2_X1 s5_U30 ( .A(randomS5[1]), .B(randomS5[9]), .Z(s5_n4) );
  XNOR2_X1 s5_U29 ( .A(s5_n2), .B(s5_n1), .ZN(s5_refreshed[24]) );
  XNOR2_X1 s5_U28 ( .A(s5_concat[24]), .B(randomS5[16]), .ZN(s5_n1) );
  XOR2_X1 s5_U27 ( .A(randomS5[0]), .B(randomS5[8]), .Z(s5_n2) );
  XOR2_X1 s5_U26 ( .A(randomS5[23]), .B(s5_concat[23]), .Z(s5_refreshed[23])
         );
  XOR2_X1 s5_U25 ( .A(randomS5[22]), .B(s5_concat[22]), .Z(s5_refreshed[22])
         );
  XOR2_X1 s5_U24 ( .A(randomS5[21]), .B(s5_concat[21]), .Z(s5_refreshed[21])
         );
  XOR2_X1 s5_U23 ( .A(randomS5[20]), .B(s5_concat[20]), .Z(s5_refreshed[20])
         );
  XOR2_X1 s5_U22 ( .A(randomS5[19]), .B(s5_concat[19]), .Z(s5_refreshed[19])
         );
  XOR2_X1 s5_U21 ( .A(randomS5[18]), .B(s5_concat[18]), .Z(s5_refreshed[18])
         );
  XOR2_X1 s5_U20 ( .A(randomS5[17]), .B(s5_concat[17]), .Z(s5_refreshed[17])
         );
  XOR2_X1 s5_U19 ( .A(randomS5[16]), .B(s5_concat[16]), .Z(s5_refreshed[16])
         );
  XOR2_X1 s5_U18 ( .A(randomS5[15]), .B(s5_concat[15]), .Z(s5_refreshed[15])
         );
  XOR2_X1 s5_U17 ( .A(randomS5[14]), .B(s5_concat[14]), .Z(s5_refreshed[14])
         );
  XOR2_X1 s5_U16 ( .A(randomS5[13]), .B(s5_concat[13]), .Z(s5_refreshed[13])
         );
  XOR2_X1 s5_U15 ( .A(randomS5[12]), .B(s5_concat[12]), .Z(s5_refreshed[12])
         );
  XOR2_X1 s5_U14 ( .A(randomS5[11]), .B(s5_concat[11]), .Z(s5_refreshed[11])
         );
  XOR2_X1 s5_U13 ( .A(randomS5[10]), .B(s5_concat[10]), .Z(s5_refreshed[10])
         );
  XOR2_X1 s5_U12 ( .A(randomS5[9]), .B(s5_concat[9]), .Z(s5_refreshed[9]) );
  XOR2_X1 s5_U11 ( .A(randomS5[8]), .B(s5_concat[8]), .Z(s5_refreshed[8]) );
  XOR2_X1 s5_U10 ( .A(randomS5[7]), .B(s5_concat[7]), .Z(s5_refreshed[7]) );
  XOR2_X1 s5_U9 ( .A(randomS5[6]), .B(s5_concat[6]), .Z(s5_refreshed[6]) );
  XOR2_X1 s5_U8 ( .A(randomS5[5]), .B(s5_concat[5]), .Z(s5_refreshed[5]) );
  XOR2_X1 s5_U7 ( .A(randomS5[4]), .B(s5_concat[4]), .Z(s5_refreshed[4]) );
  XOR2_X1 s5_U6 ( .A(randomS5[3]), .B(s5_concat[3]), .Z(s5_refreshed[3]) );
  XOR2_X1 s5_U5 ( .A(randomS5[2]), .B(s5_concat[2]), .Z(s5_refreshed[2]) );
  XOR2_X1 s5_U4 ( .A(randomS5[1]), .B(s5_concat[1]), .Z(s5_refreshed[1]) );
  XOR2_X1 s5_U3 ( .A(randomS5[0]), .B(s5_concat[0]), .Z(s5_refreshed[0]) );
  DFF_X1 s5_regOut_reg_0__0__0_ ( .D(s5_refreshed[0]), .CK(clk), .Q(
        s5_regOut[0]), .QN() );
  DFF_X1 s5_regOut_reg_0__0__1_ ( .D(s5_refreshed[1]), .CK(clk), .Q(
        s5_regOut[1]), .QN() );
  DFF_X1 s5_regOut_reg_0__0__2_ ( .D(s5_refreshed[2]), .CK(clk), .Q(
        s5_regOut[2]), .QN() );
  DFF_X1 s5_regOut_reg_0__0__3_ ( .D(s5_refreshed[3]), .CK(clk), .Q(
        s5_regOut[3]), .QN() );
  DFF_X1 s5_regOut_reg_0__0__4_ ( .D(s5_refreshed[4]), .CK(clk), .Q(
        s5_regOut[4]), .QN() );
  DFF_X1 s5_regOut_reg_0__0__5_ ( .D(s5_refreshed[5]), .CK(clk), .Q(
        s5_regOut[5]), .QN() );
  DFF_X1 s5_regOut_reg_0__0__6_ ( .D(s5_refreshed[6]), .CK(clk), .Q(
        s5_regOut[6]), .QN() );
  DFF_X1 s5_regOut_reg_0__0__7_ ( .D(s5_refreshed[7]), .CK(clk), .Q(
        s5_regOut[7]), .QN() );
  DFF_X1 s5_regOut_reg_0__1__0_ ( .D(s5_refreshed[8]), .CK(clk), .Q(
        s5_regOut[8]), .QN() );
  DFF_X1 s5_regOut_reg_0__1__1_ ( .D(s5_refreshed[9]), .CK(clk), .Q(
        s5_regOut[9]), .QN() );
  DFF_X1 s5_regOut_reg_0__1__2_ ( .D(s5_refreshed[10]), .CK(clk), .Q(
        s5_regOut[10]), .QN() );
  DFF_X1 s5_regOut_reg_0__1__3_ ( .D(s5_refreshed[11]), .CK(clk), .Q(
        s5_regOut[11]), .QN() );
  DFF_X1 s5_regOut_reg_0__1__4_ ( .D(s5_refreshed[12]), .CK(clk), .Q(
        s5_regOut[12]), .QN() );
  DFF_X1 s5_regOut_reg_0__1__5_ ( .D(s5_refreshed[13]), .CK(clk), .Q(
        s5_regOut[13]), .QN() );
  DFF_X1 s5_regOut_reg_0__1__6_ ( .D(s5_refreshed[14]), .CK(clk), .Q(
        s5_regOut[14]), .QN() );
  DFF_X1 s5_regOut_reg_0__1__7_ ( .D(s5_refreshed[15]), .CK(clk), .Q(
        s5_regOut[15]), .QN() );
  DFF_X1 s5_regOut_reg_1__0__0_ ( .D(s5_refreshed[16]), .CK(clk), .Q(
        s5_regOut[16]), .QN() );
  DFF_X1 s5_regOut_reg_1__0__1_ ( .D(s5_refreshed[17]), .CK(clk), .Q(
        s5_regOut[17]), .QN() );
  DFF_X1 s5_regOut_reg_1__0__2_ ( .D(s5_refreshed[18]), .CK(clk), .Q(
        s5_regOut[18]), .QN() );
  DFF_X1 s5_regOut_reg_1__0__3_ ( .D(s5_refreshed[19]), .CK(clk), .Q(
        s5_regOut[19]), .QN() );
  DFF_X1 s5_regOut_reg_1__0__4_ ( .D(s5_refreshed[20]), .CK(clk), .Q(
        s5_regOut[20]), .QN() );
  DFF_X1 s5_regOut_reg_1__0__5_ ( .D(s5_refreshed[21]), .CK(clk), .Q(
        s5_regOut[21]), .QN() );
  DFF_X1 s5_regOut_reg_1__0__6_ ( .D(s5_refreshed[22]), .CK(clk), .Q(
        s5_regOut[22]), .QN() );
  DFF_X1 s5_regOut_reg_1__0__7_ ( .D(s5_refreshed[23]), .CK(clk), .Q(
        s5_regOut[23]), .QN() );
  DFF_X1 s5_regOut_reg_1__1__0_ ( .D(s5_refreshed[24]), .CK(clk), .Q(
        s5_regOut[24]), .QN() );
  DFF_X1 s5_regOut_reg_1__1__1_ ( .D(s5_refreshed[25]), .CK(clk), .Q(
        s5_regOut[25]), .QN() );
  DFF_X1 s5_regOut_reg_1__1__2_ ( .D(s5_refreshed[26]), .CK(clk), .Q(
        s5_regOut[26]), .QN() );
  DFF_X1 s5_regOut_reg_1__1__3_ ( .D(s5_refreshed[27]), .CK(clk), .Q(
        s5_regOut[27]), .QN() );
  DFF_X1 s5_regOut_reg_1__1__4_ ( .D(s5_refreshed[28]), .CK(clk), .Q(
        s5_regOut[28]), .QN() );
  DFF_X1 s5_regOut_reg_1__1__5_ ( .D(s5_refreshed[29]), .CK(clk), .Q(
        s5_regOut[29]), .QN() );
  DFF_X1 s5_regOut_reg_1__1__6_ ( .D(s5_refreshed[30]), .CK(clk), .Q(
        s5_regOut[30]), .QN() );
  DFF_X1 s5_regOut_reg_1__1__7_ ( .D(s5_refreshed[31]), .CK(clk), .Q(
        s5_regOut[31]), .QN() );
  XNOR2_X1 s5_mul1_1_1_U29 ( .A(s5_mul1_1_1_n77), .B(s5_mul1_1_1_n76), .ZN(
        s5_concat[27]) );
  NAND2_X1 s5_mul1_1_1_U28 ( .A1(stage4Out[23]), .A2(stage4Out[19]), .ZN(
        s5_mul1_1_1_n76) );
  XOR2_X1 s5_mul1_1_1_U27 ( .A(s5_mul1_1_1_n75), .B(s5_mul1_1_1_n74), .Z(
        s5_mul1_1_1_n77) );
  XNOR2_X1 s5_mul1_1_1_U26 ( .A(s5_mul1_1_1_n73), .B(s5_mul1_1_1_n72), .ZN(
        s5_concat[26]) );
  NAND2_X1 s5_mul1_1_1_U25 ( .A1(stage4Out[22]), .A2(stage4Out[18]), .ZN(
        s5_mul1_1_1_n72) );
  XOR2_X1 s5_mul1_1_1_U24 ( .A(s5_mul1_1_1_n74), .B(s5_mul1_1_1_n71), .Z(
        s5_mul1_1_1_n73) );
  NOR2_X1 s5_mul1_1_1_U23 ( .A1(s5_mul1_1_1_n70), .A2(s5_mul1_1_1_n69), .ZN(
        s5_mul1_1_1_n74) );
  XNOR2_X1 s5_mul1_1_1_U22 ( .A(stage4Out[22]), .B(stage4Out[23]), .ZN(
        s5_mul1_1_1_n69) );
  XNOR2_X1 s5_mul1_1_1_U21 ( .A(stage4Out[18]), .B(stage4Out[19]), .ZN(
        s5_mul1_1_1_n70) );
  XNOR2_X1 s5_mul1_1_1_U20 ( .A(s5_mul1_1_1_n68), .B(s5_mul1_1_1_n67), .ZN(
        s5_concat[25]) );
  NAND2_X1 s5_mul1_1_1_U19 ( .A1(stage4Out[21]), .A2(stage4Out[17]), .ZN(
        s5_mul1_1_1_n67) );
  XOR2_X1 s5_mul1_1_1_U18 ( .A(s5_mul1_1_1_n75), .B(s5_mul1_1_1_n66), .Z(
        s5_mul1_1_1_n68) );
  XNOR2_X1 s5_mul1_1_1_U17 ( .A(s5_mul1_1_1_n65), .B(s5_mul1_1_1_n64), .ZN(
        s5_mul1_1_1_n75) );
  NAND2_X1 s5_mul1_1_1_U16 ( .A1(s5_mul1_1_1_n63), .A2(s5_mul1_1_1_n62), .ZN(
        s5_mul1_1_1_n64) );
  XNOR2_X1 s5_mul1_1_1_U15 ( .A(s5_mul1_1_1_n61), .B(s5_mul1_1_1_n60), .ZN(
        s5_mul1_1_1_n62) );
  XNOR2_X1 s5_mul1_1_1_U14 ( .A(s5_mul1_1_1_n59), .B(s5_mul1_1_1_n58), .ZN(
        s5_mul1_1_1_n63) );
  XNOR2_X1 s5_mul1_1_1_U13 ( .A(s5_mul1_1_1_n57), .B(s5_mul1_1_1_n56), .ZN(
        s5_concat[24]) );
  NAND2_X1 s5_mul1_1_1_U12 ( .A1(stage4Out[20]), .A2(stage4Out[16]), .ZN(
        s5_mul1_1_1_n56) );
  XOR2_X1 s5_mul1_1_1_U11 ( .A(s5_mul1_1_1_n66), .B(s5_mul1_1_1_n71), .Z(
        s5_mul1_1_1_n57) );
  XNOR2_X1 s5_mul1_1_1_U10 ( .A(s5_mul1_1_1_n55), .B(s5_mul1_1_1_n65), .ZN(
        s5_mul1_1_1_n71) );
  NOR2_X1 s5_mul1_1_1_U9 ( .A1(s5_mul1_1_1_n61), .A2(s5_mul1_1_1_n59), .ZN(
        s5_mul1_1_1_n65) );
  XNOR2_X1 s5_mul1_1_1_U8 ( .A(stage4Out[20]), .B(stage4Out[22]), .ZN(
        s5_mul1_1_1_n59) );
  XNOR2_X1 s5_mul1_1_1_U7 ( .A(stage4Out[16]), .B(stage4Out[18]), .ZN(
        s5_mul1_1_1_n61) );
  NAND2_X1 s5_mul1_1_1_U6 ( .A1(s5_mul1_1_1_n58), .A2(s5_mul1_1_1_n60), .ZN(
        s5_mul1_1_1_n55) );
  XOR2_X1 s5_mul1_1_1_U5 ( .A(stage4Out[17]), .B(stage4Out[19]), .Z(
        s5_mul1_1_1_n60) );
  XOR2_X1 s5_mul1_1_1_U4 ( .A(stage4Out[21]), .B(stage4Out[23]), .Z(
        s5_mul1_1_1_n58) );
  NOR2_X1 s5_mul1_1_1_U3 ( .A1(s5_mul1_1_1_n54), .A2(s5_mul1_1_1_n53), .ZN(
        s5_mul1_1_1_n66) );
  XNOR2_X1 s5_mul1_1_1_U2 ( .A(stage4Out[20]), .B(stage4Out[21]), .ZN(
        s5_mul1_1_1_n53) );
  XNOR2_X1 s5_mul1_1_1_U1 ( .A(stage4Out[16]), .B(stage4Out[17]), .ZN(
        s5_mul1_1_1_n54) );
  XNOR2_X1 s5_mul1_1_0_U29 ( .A(s5_mul1_1_0_n77), .B(s5_mul1_1_0_n76), .ZN(
        s5_concat[19]) );
  NAND2_X1 s5_mul1_1_0_U28 ( .A1(stage4Out[23]), .A2(stage4Out[7]), .ZN(
        s5_mul1_1_0_n76) );
  XOR2_X1 s5_mul1_1_0_U27 ( .A(s5_mul1_1_0_n75), .B(s5_mul1_1_0_n74), .Z(
        s5_mul1_1_0_n77) );
  XNOR2_X1 s5_mul1_1_0_U26 ( .A(s5_mul1_1_0_n73), .B(s5_mul1_1_0_n72), .ZN(
        s5_concat[18]) );
  NAND2_X1 s5_mul1_1_0_U25 ( .A1(stage4Out[22]), .A2(stage4Out[6]), .ZN(
        s5_mul1_1_0_n72) );
  XOR2_X1 s5_mul1_1_0_U24 ( .A(s5_mul1_1_0_n74), .B(s5_mul1_1_0_n71), .Z(
        s5_mul1_1_0_n73) );
  NOR2_X1 s5_mul1_1_0_U23 ( .A1(s5_mul1_1_0_n70), .A2(s5_mul1_1_0_n69), .ZN(
        s5_mul1_1_0_n74) );
  XNOR2_X1 s5_mul1_1_0_U22 ( .A(stage4Out[22]), .B(stage4Out[23]), .ZN(
        s5_mul1_1_0_n69) );
  XNOR2_X1 s5_mul1_1_0_U21 ( .A(stage4Out[6]), .B(stage4Out[7]), .ZN(
        s5_mul1_1_0_n70) );
  XNOR2_X1 s5_mul1_1_0_U20 ( .A(s5_mul1_1_0_n68), .B(s5_mul1_1_0_n67), .ZN(
        s5_concat[17]) );
  NAND2_X1 s5_mul1_1_0_U19 ( .A1(stage4Out[21]), .A2(stage4Out[5]), .ZN(
        s5_mul1_1_0_n67) );
  XOR2_X1 s5_mul1_1_0_U18 ( .A(s5_mul1_1_0_n75), .B(s5_mul1_1_0_n66), .Z(
        s5_mul1_1_0_n68) );
  XNOR2_X1 s5_mul1_1_0_U17 ( .A(s5_mul1_1_0_n65), .B(s5_mul1_1_0_n64), .ZN(
        s5_mul1_1_0_n75) );
  NAND2_X1 s5_mul1_1_0_U16 ( .A1(s5_mul1_1_0_n63), .A2(s5_mul1_1_0_n62), .ZN(
        s5_mul1_1_0_n64) );
  XNOR2_X1 s5_mul1_1_0_U15 ( .A(s5_mul1_1_0_n61), .B(s5_mul1_1_0_n60), .ZN(
        s5_mul1_1_0_n62) );
  XNOR2_X1 s5_mul1_1_0_U14 ( .A(s5_mul1_1_0_n59), .B(s5_mul1_1_0_n58), .ZN(
        s5_mul1_1_0_n63) );
  XNOR2_X1 s5_mul1_1_0_U13 ( .A(s5_mul1_1_0_n57), .B(s5_mul1_1_0_n56), .ZN(
        s5_concat[16]) );
  NAND2_X1 s5_mul1_1_0_U12 ( .A1(stage4Out[20]), .A2(stage4Out[4]), .ZN(
        s5_mul1_1_0_n56) );
  XOR2_X1 s5_mul1_1_0_U11 ( .A(s5_mul1_1_0_n66), .B(s5_mul1_1_0_n71), .Z(
        s5_mul1_1_0_n57) );
  XNOR2_X1 s5_mul1_1_0_U10 ( .A(s5_mul1_1_0_n55), .B(s5_mul1_1_0_n65), .ZN(
        s5_mul1_1_0_n71) );
  NOR2_X1 s5_mul1_1_0_U9 ( .A1(s5_mul1_1_0_n61), .A2(s5_mul1_1_0_n59), .ZN(
        s5_mul1_1_0_n65) );
  XNOR2_X1 s5_mul1_1_0_U8 ( .A(stage4Out[20]), .B(stage4Out[22]), .ZN(
        s5_mul1_1_0_n59) );
  XNOR2_X1 s5_mul1_1_0_U7 ( .A(stage4Out[4]), .B(stage4Out[6]), .ZN(
        s5_mul1_1_0_n61) );
  NAND2_X1 s5_mul1_1_0_U6 ( .A1(s5_mul1_1_0_n58), .A2(s5_mul1_1_0_n60), .ZN(
        s5_mul1_1_0_n55) );
  XOR2_X1 s5_mul1_1_0_U5 ( .A(stage4Out[5]), .B(stage4Out[7]), .Z(
        s5_mul1_1_0_n60) );
  XOR2_X1 s5_mul1_1_0_U4 ( .A(stage4Out[21]), .B(stage4Out[23]), .Z(
        s5_mul1_1_0_n58) );
  NOR2_X1 s5_mul1_1_0_U3 ( .A1(s5_mul1_1_0_n54), .A2(s5_mul1_1_0_n53), .ZN(
        s5_mul1_1_0_n66) );
  XNOR2_X1 s5_mul1_1_0_U2 ( .A(stage4Out[20]), .B(stage4Out[21]), .ZN(
        s5_mul1_1_0_n53) );
  XNOR2_X1 s5_mul1_1_0_U1 ( .A(stage4Out[4]), .B(stage4Out[5]), .ZN(
        s5_mul1_1_0_n54) );
  XNOR2_X1 s5_mul1_0_1_U29 ( .A(s5_mul1_0_1_n77), .B(s5_mul1_0_1_n76), .ZN(
        s5_concat[11]) );
  NAND2_X1 s5_mul1_0_1_U28 ( .A1(stage4Out[11]), .A2(stage4Out[19]), .ZN(
        s5_mul1_0_1_n76) );
  XOR2_X1 s5_mul1_0_1_U27 ( .A(s5_mul1_0_1_n75), .B(s5_mul1_0_1_n74), .Z(
        s5_mul1_0_1_n77) );
  XNOR2_X1 s5_mul1_0_1_U26 ( .A(s5_mul1_0_1_n73), .B(s5_mul1_0_1_n72), .ZN(
        s5_concat[10]) );
  NAND2_X1 s5_mul1_0_1_U25 ( .A1(stage4Out[10]), .A2(stage4Out[18]), .ZN(
        s5_mul1_0_1_n72) );
  XOR2_X1 s5_mul1_0_1_U24 ( .A(s5_mul1_0_1_n74), .B(s5_mul1_0_1_n71), .Z(
        s5_mul1_0_1_n73) );
  NOR2_X1 s5_mul1_0_1_U23 ( .A1(s5_mul1_0_1_n70), .A2(s5_mul1_0_1_n69), .ZN(
        s5_mul1_0_1_n74) );
  XNOR2_X1 s5_mul1_0_1_U22 ( .A(stage4Out[10]), .B(stage4Out[11]), .ZN(
        s5_mul1_0_1_n69) );
  XNOR2_X1 s5_mul1_0_1_U21 ( .A(stage4Out[18]), .B(stage4Out[19]), .ZN(
        s5_mul1_0_1_n70) );
  XNOR2_X1 s5_mul1_0_1_U20 ( .A(s5_mul1_0_1_n68), .B(s5_mul1_0_1_n67), .ZN(
        s5_concat[9]) );
  NAND2_X1 s5_mul1_0_1_U19 ( .A1(stage4Out[9]), .A2(stage4Out[17]), .ZN(
        s5_mul1_0_1_n67) );
  XOR2_X1 s5_mul1_0_1_U18 ( .A(s5_mul1_0_1_n75), .B(s5_mul1_0_1_n66), .Z(
        s5_mul1_0_1_n68) );
  XNOR2_X1 s5_mul1_0_1_U17 ( .A(s5_mul1_0_1_n65), .B(s5_mul1_0_1_n64), .ZN(
        s5_mul1_0_1_n75) );
  NAND2_X1 s5_mul1_0_1_U16 ( .A1(s5_mul1_0_1_n63), .A2(s5_mul1_0_1_n62), .ZN(
        s5_mul1_0_1_n64) );
  XNOR2_X1 s5_mul1_0_1_U15 ( .A(s5_mul1_0_1_n61), .B(s5_mul1_0_1_n60), .ZN(
        s5_mul1_0_1_n62) );
  XNOR2_X1 s5_mul1_0_1_U14 ( .A(s5_mul1_0_1_n59), .B(s5_mul1_0_1_n58), .ZN(
        s5_mul1_0_1_n63) );
  XNOR2_X1 s5_mul1_0_1_U13 ( .A(s5_mul1_0_1_n57), .B(s5_mul1_0_1_n56), .ZN(
        s5_concat[8]) );
  NAND2_X1 s5_mul1_0_1_U12 ( .A1(stage4Out[8]), .A2(stage4Out[16]), .ZN(
        s5_mul1_0_1_n56) );
  XOR2_X1 s5_mul1_0_1_U11 ( .A(s5_mul1_0_1_n66), .B(s5_mul1_0_1_n71), .Z(
        s5_mul1_0_1_n57) );
  XNOR2_X1 s5_mul1_0_1_U10 ( .A(s5_mul1_0_1_n55), .B(s5_mul1_0_1_n65), .ZN(
        s5_mul1_0_1_n71) );
  NOR2_X1 s5_mul1_0_1_U9 ( .A1(s5_mul1_0_1_n61), .A2(s5_mul1_0_1_n59), .ZN(
        s5_mul1_0_1_n65) );
  XNOR2_X1 s5_mul1_0_1_U8 ( .A(stage4Out[8]), .B(stage4Out[10]), .ZN(
        s5_mul1_0_1_n59) );
  XNOR2_X1 s5_mul1_0_1_U7 ( .A(stage4Out[16]), .B(stage4Out[18]), .ZN(
        s5_mul1_0_1_n61) );
  NAND2_X1 s5_mul1_0_1_U6 ( .A1(s5_mul1_0_1_n58), .A2(s5_mul1_0_1_n60), .ZN(
        s5_mul1_0_1_n55) );
  XOR2_X1 s5_mul1_0_1_U5 ( .A(stage4Out[17]), .B(stage4Out[19]), .Z(
        s5_mul1_0_1_n60) );
  XOR2_X1 s5_mul1_0_1_U4 ( .A(stage4Out[9]), .B(stage4Out[11]), .Z(
        s5_mul1_0_1_n58) );
  NOR2_X1 s5_mul1_0_1_U3 ( .A1(s5_mul1_0_1_n54), .A2(s5_mul1_0_1_n53), .ZN(
        s5_mul1_0_1_n66) );
  XNOR2_X1 s5_mul1_0_1_U2 ( .A(stage4Out[8]), .B(stage4Out[9]), .ZN(
        s5_mul1_0_1_n53) );
  XNOR2_X1 s5_mul1_0_1_U1 ( .A(stage4Out[16]), .B(stage4Out[17]), .ZN(
        s5_mul1_0_1_n54) );
  XNOR2_X1 s5_mul1_0_0_U29 ( .A(s5_mul1_0_0_n77), .B(s5_mul1_0_0_n76), .ZN(
        s5_concat[3]) );
  NAND2_X1 s5_mul1_0_0_U28 ( .A1(stage4Out[11]), .A2(stage4Out[7]), .ZN(
        s5_mul1_0_0_n76) );
  XOR2_X1 s5_mul1_0_0_U27 ( .A(s5_mul1_0_0_n75), .B(s5_mul1_0_0_n74), .Z(
        s5_mul1_0_0_n77) );
  XNOR2_X1 s5_mul1_0_0_U26 ( .A(s5_mul1_0_0_n73), .B(s5_mul1_0_0_n72), .ZN(
        s5_concat[2]) );
  NAND2_X1 s5_mul1_0_0_U25 ( .A1(stage4Out[10]), .A2(stage4Out[6]), .ZN(
        s5_mul1_0_0_n72) );
  XOR2_X1 s5_mul1_0_0_U24 ( .A(s5_mul1_0_0_n74), .B(s5_mul1_0_0_n71), .Z(
        s5_mul1_0_0_n73) );
  NOR2_X1 s5_mul1_0_0_U23 ( .A1(s5_mul1_0_0_n70), .A2(s5_mul1_0_0_n69), .ZN(
        s5_mul1_0_0_n74) );
  XNOR2_X1 s5_mul1_0_0_U22 ( .A(stage4Out[10]), .B(stage4Out[11]), .ZN(
        s5_mul1_0_0_n69) );
  XNOR2_X1 s5_mul1_0_0_U21 ( .A(stage4Out[6]), .B(stage4Out[7]), .ZN(
        s5_mul1_0_0_n70) );
  XNOR2_X1 s5_mul1_0_0_U20 ( .A(s5_mul1_0_0_n68), .B(s5_mul1_0_0_n67), .ZN(
        s5_concat[1]) );
  NAND2_X1 s5_mul1_0_0_U19 ( .A1(stage4Out[9]), .A2(stage4Out[5]), .ZN(
        s5_mul1_0_0_n67) );
  XOR2_X1 s5_mul1_0_0_U18 ( .A(s5_mul1_0_0_n75), .B(s5_mul1_0_0_n66), .Z(
        s5_mul1_0_0_n68) );
  XNOR2_X1 s5_mul1_0_0_U17 ( .A(s5_mul1_0_0_n65), .B(s5_mul1_0_0_n64), .ZN(
        s5_mul1_0_0_n75) );
  NAND2_X1 s5_mul1_0_0_U16 ( .A1(s5_mul1_0_0_n63), .A2(s5_mul1_0_0_n62), .ZN(
        s5_mul1_0_0_n64) );
  XNOR2_X1 s5_mul1_0_0_U15 ( .A(s5_mul1_0_0_n61), .B(s5_mul1_0_0_n60), .ZN(
        s5_mul1_0_0_n62) );
  XNOR2_X1 s5_mul1_0_0_U14 ( .A(s5_mul1_0_0_n59), .B(s5_mul1_0_0_n58), .ZN(
        s5_mul1_0_0_n63) );
  XNOR2_X1 s5_mul1_0_0_U13 ( .A(s5_mul1_0_0_n57), .B(s5_mul1_0_0_n56), .ZN(
        s5_concat[0]) );
  NAND2_X1 s5_mul1_0_0_U12 ( .A1(stage4Out[8]), .A2(stage4Out[4]), .ZN(
        s5_mul1_0_0_n56) );
  XOR2_X1 s5_mul1_0_0_U11 ( .A(s5_mul1_0_0_n66), .B(s5_mul1_0_0_n71), .Z(
        s5_mul1_0_0_n57) );
  XNOR2_X1 s5_mul1_0_0_U10 ( .A(s5_mul1_0_0_n55), .B(s5_mul1_0_0_n65), .ZN(
        s5_mul1_0_0_n71) );
  NOR2_X1 s5_mul1_0_0_U9 ( .A1(s5_mul1_0_0_n61), .A2(s5_mul1_0_0_n59), .ZN(
        s5_mul1_0_0_n65) );
  XNOR2_X1 s5_mul1_0_0_U8 ( .A(stage4Out[8]), .B(stage4Out[10]), .ZN(
        s5_mul1_0_0_n59) );
  XNOR2_X1 s5_mul1_0_0_U7 ( .A(stage4Out[4]), .B(stage4Out[6]), .ZN(
        s5_mul1_0_0_n61) );
  NAND2_X1 s5_mul1_0_0_U6 ( .A1(s5_mul1_0_0_n58), .A2(s5_mul1_0_0_n60), .ZN(
        s5_mul1_0_0_n55) );
  XOR2_X1 s5_mul1_0_0_U5 ( .A(stage4Out[5]), .B(stage4Out[7]), .Z(
        s5_mul1_0_0_n60) );
  XOR2_X1 s5_mul1_0_0_U4 ( .A(stage4Out[9]), .B(stage4Out[11]), .Z(
        s5_mul1_0_0_n58) );
  NOR2_X1 s5_mul1_0_0_U3 ( .A1(s5_mul1_0_0_n54), .A2(s5_mul1_0_0_n53), .ZN(
        s5_mul1_0_0_n66) );
  XNOR2_X1 s5_mul1_0_0_U2 ( .A(stage4Out[8]), .B(stage4Out[9]), .ZN(
        s5_mul1_0_0_n53) );
  XNOR2_X1 s5_mul1_0_0_U1 ( .A(stage4Out[4]), .B(stage4Out[5]), .ZN(
        s5_mul1_0_0_n54) );
  XNOR2_X1 s5_mul2_1_1_U29 ( .A(s5_mul2_1_1_n77), .B(s5_mul2_1_1_n76), .ZN(
        s5_concat[31]) );
  NAND2_X1 s5_mul2_1_1_U28 ( .A1(stage4Out[19]), .A2(stage4Out[15]), .ZN(
        s5_mul2_1_1_n76) );
  XOR2_X1 s5_mul2_1_1_U27 ( .A(s5_mul2_1_1_n75), .B(s5_mul2_1_1_n74), .Z(
        s5_mul2_1_1_n77) );
  XNOR2_X1 s5_mul2_1_1_U26 ( .A(s5_mul2_1_1_n73), .B(s5_mul2_1_1_n72), .ZN(
        s5_concat[30]) );
  NAND2_X1 s5_mul2_1_1_U25 ( .A1(stage4Out[18]), .A2(stage4Out[14]), .ZN(
        s5_mul2_1_1_n72) );
  XOR2_X1 s5_mul2_1_1_U24 ( .A(s5_mul2_1_1_n74), .B(s5_mul2_1_1_n71), .Z(
        s5_mul2_1_1_n73) );
  NOR2_X1 s5_mul2_1_1_U23 ( .A1(s5_mul2_1_1_n70), .A2(s5_mul2_1_1_n69), .ZN(
        s5_mul2_1_1_n74) );
  XNOR2_X1 s5_mul2_1_1_U22 ( .A(stage4Out[18]), .B(stage4Out[19]), .ZN(
        s5_mul2_1_1_n69) );
  XNOR2_X1 s5_mul2_1_1_U21 ( .A(stage4Out[14]), .B(stage4Out[15]), .ZN(
        s5_mul2_1_1_n70) );
  XNOR2_X1 s5_mul2_1_1_U20 ( .A(s5_mul2_1_1_n68), .B(s5_mul2_1_1_n67), .ZN(
        s5_concat[29]) );
  NAND2_X1 s5_mul2_1_1_U19 ( .A1(stage4Out[17]), .A2(stage4Out[13]), .ZN(
        s5_mul2_1_1_n67) );
  XOR2_X1 s5_mul2_1_1_U18 ( .A(s5_mul2_1_1_n75), .B(s5_mul2_1_1_n66), .Z(
        s5_mul2_1_1_n68) );
  XNOR2_X1 s5_mul2_1_1_U17 ( .A(s5_mul2_1_1_n65), .B(s5_mul2_1_1_n64), .ZN(
        s5_mul2_1_1_n75) );
  NAND2_X1 s5_mul2_1_1_U16 ( .A1(s5_mul2_1_1_n63), .A2(s5_mul2_1_1_n62), .ZN(
        s5_mul2_1_1_n64) );
  XNOR2_X1 s5_mul2_1_1_U15 ( .A(s5_mul2_1_1_n61), .B(s5_mul2_1_1_n60), .ZN(
        s5_mul2_1_1_n62) );
  XNOR2_X1 s5_mul2_1_1_U14 ( .A(s5_mul2_1_1_n59), .B(s5_mul2_1_1_n58), .ZN(
        s5_mul2_1_1_n63) );
  XNOR2_X1 s5_mul2_1_1_U13 ( .A(s5_mul2_1_1_n57), .B(s5_mul2_1_1_n56), .ZN(
        s5_concat[28]) );
  NAND2_X1 s5_mul2_1_1_U12 ( .A1(stage4Out[16]), .A2(stage4Out[12]), .ZN(
        s5_mul2_1_1_n56) );
  XOR2_X1 s5_mul2_1_1_U11 ( .A(s5_mul2_1_1_n66), .B(s5_mul2_1_1_n71), .Z(
        s5_mul2_1_1_n57) );
  XNOR2_X1 s5_mul2_1_1_U10 ( .A(s5_mul2_1_1_n55), .B(s5_mul2_1_1_n65), .ZN(
        s5_mul2_1_1_n71) );
  NOR2_X1 s5_mul2_1_1_U9 ( .A1(s5_mul2_1_1_n61), .A2(s5_mul2_1_1_n59), .ZN(
        s5_mul2_1_1_n65) );
  XNOR2_X1 s5_mul2_1_1_U8 ( .A(stage4Out[16]), .B(stage4Out[18]), .ZN(
        s5_mul2_1_1_n59) );
  XNOR2_X1 s5_mul2_1_1_U7 ( .A(stage4Out[12]), .B(stage4Out[14]), .ZN(
        s5_mul2_1_1_n61) );
  NAND2_X1 s5_mul2_1_1_U6 ( .A1(s5_mul2_1_1_n58), .A2(s5_mul2_1_1_n60), .ZN(
        s5_mul2_1_1_n55) );
  XOR2_X1 s5_mul2_1_1_U5 ( .A(stage4Out[13]), .B(stage4Out[15]), .Z(
        s5_mul2_1_1_n60) );
  XOR2_X1 s5_mul2_1_1_U4 ( .A(stage4Out[17]), .B(stage4Out[19]), .Z(
        s5_mul2_1_1_n58) );
  NOR2_X1 s5_mul2_1_1_U3 ( .A1(s5_mul2_1_1_n54), .A2(s5_mul2_1_1_n53), .ZN(
        s5_mul2_1_1_n66) );
  XNOR2_X1 s5_mul2_1_1_U2 ( .A(stage4Out[16]), .B(stage4Out[17]), .ZN(
        s5_mul2_1_1_n53) );
  XNOR2_X1 s5_mul2_1_1_U1 ( .A(stage4Out[12]), .B(stage4Out[13]), .ZN(
        s5_mul2_1_1_n54) );
  XNOR2_X1 s5_mul2_1_0_U29 ( .A(s5_mul2_1_0_n77), .B(s5_mul2_1_0_n76), .ZN(
        s5_concat[23]) );
  NAND2_X1 s5_mul2_1_0_U28 ( .A1(stage4Out[19]), .A2(stage4Out[3]), .ZN(
        s5_mul2_1_0_n76) );
  XOR2_X1 s5_mul2_1_0_U27 ( .A(s5_mul2_1_0_n75), .B(s5_mul2_1_0_n74), .Z(
        s5_mul2_1_0_n77) );
  XNOR2_X1 s5_mul2_1_0_U26 ( .A(s5_mul2_1_0_n73), .B(s5_mul2_1_0_n72), .ZN(
        s5_concat[22]) );
  NAND2_X1 s5_mul2_1_0_U25 ( .A1(stage4Out[18]), .A2(stage4Out[2]), .ZN(
        s5_mul2_1_0_n72) );
  XOR2_X1 s5_mul2_1_0_U24 ( .A(s5_mul2_1_0_n74), .B(s5_mul2_1_0_n71), .Z(
        s5_mul2_1_0_n73) );
  NOR2_X1 s5_mul2_1_0_U23 ( .A1(s5_mul2_1_0_n70), .A2(s5_mul2_1_0_n69), .ZN(
        s5_mul2_1_0_n74) );
  XNOR2_X1 s5_mul2_1_0_U22 ( .A(stage4Out[18]), .B(stage4Out[19]), .ZN(
        s5_mul2_1_0_n69) );
  XNOR2_X1 s5_mul2_1_0_U21 ( .A(stage4Out[2]), .B(stage4Out[3]), .ZN(
        s5_mul2_1_0_n70) );
  XNOR2_X1 s5_mul2_1_0_U20 ( .A(s5_mul2_1_0_n68), .B(s5_mul2_1_0_n67), .ZN(
        s5_concat[21]) );
  NAND2_X1 s5_mul2_1_0_U19 ( .A1(stage4Out[17]), .A2(stage4Out[1]), .ZN(
        s5_mul2_1_0_n67) );
  XOR2_X1 s5_mul2_1_0_U18 ( .A(s5_mul2_1_0_n75), .B(s5_mul2_1_0_n66), .Z(
        s5_mul2_1_0_n68) );
  XNOR2_X1 s5_mul2_1_0_U17 ( .A(s5_mul2_1_0_n65), .B(s5_mul2_1_0_n64), .ZN(
        s5_mul2_1_0_n75) );
  NAND2_X1 s5_mul2_1_0_U16 ( .A1(s5_mul2_1_0_n63), .A2(s5_mul2_1_0_n62), .ZN(
        s5_mul2_1_0_n64) );
  XNOR2_X1 s5_mul2_1_0_U15 ( .A(s5_mul2_1_0_n61), .B(s5_mul2_1_0_n60), .ZN(
        s5_mul2_1_0_n62) );
  XNOR2_X1 s5_mul2_1_0_U14 ( .A(s5_mul2_1_0_n59), .B(s5_mul2_1_0_n58), .ZN(
        s5_mul2_1_0_n63) );
  XNOR2_X1 s5_mul2_1_0_U13 ( .A(s5_mul2_1_0_n57), .B(s5_mul2_1_0_n56), .ZN(
        s5_concat[20]) );
  NAND2_X1 s5_mul2_1_0_U12 ( .A1(stage4Out[16]), .A2(stage4Out[0]), .ZN(
        s5_mul2_1_0_n56) );
  XOR2_X1 s5_mul2_1_0_U11 ( .A(s5_mul2_1_0_n66), .B(s5_mul2_1_0_n71), .Z(
        s5_mul2_1_0_n57) );
  XNOR2_X1 s5_mul2_1_0_U10 ( .A(s5_mul2_1_0_n55), .B(s5_mul2_1_0_n65), .ZN(
        s5_mul2_1_0_n71) );
  NOR2_X1 s5_mul2_1_0_U9 ( .A1(s5_mul2_1_0_n61), .A2(s5_mul2_1_0_n59), .ZN(
        s5_mul2_1_0_n65) );
  XNOR2_X1 s5_mul2_1_0_U8 ( .A(stage4Out[16]), .B(stage4Out[18]), .ZN(
        s5_mul2_1_0_n59) );
  XNOR2_X1 s5_mul2_1_0_U7 ( .A(stage4Out[0]), .B(stage4Out[2]), .ZN(
        s5_mul2_1_0_n61) );
  NAND2_X1 s5_mul2_1_0_U6 ( .A1(s5_mul2_1_0_n58), .A2(s5_mul2_1_0_n60), .ZN(
        s5_mul2_1_0_n55) );
  XOR2_X1 s5_mul2_1_0_U5 ( .A(stage4Out[1]), .B(stage4Out[3]), .Z(
        s5_mul2_1_0_n60) );
  XOR2_X1 s5_mul2_1_0_U4 ( .A(stage4Out[17]), .B(stage4Out[19]), .Z(
        s5_mul2_1_0_n58) );
  NOR2_X1 s5_mul2_1_0_U3 ( .A1(s5_mul2_1_0_n54), .A2(s5_mul2_1_0_n53), .ZN(
        s5_mul2_1_0_n66) );
  XNOR2_X1 s5_mul2_1_0_U2 ( .A(stage4Out[16]), .B(stage4Out[17]), .ZN(
        s5_mul2_1_0_n53) );
  XNOR2_X1 s5_mul2_1_0_U1 ( .A(stage4Out[0]), .B(stage4Out[1]), .ZN(
        s5_mul2_1_0_n54) );
  XNOR2_X1 s5_mul2_0_1_U29 ( .A(s5_mul2_0_1_n77), .B(s5_mul2_0_1_n76), .ZN(
        s5_concat[15]) );
  NAND2_X1 s5_mul2_0_1_U28 ( .A1(stage4Out[7]), .A2(stage4Out[15]), .ZN(
        s5_mul2_0_1_n76) );
  XOR2_X1 s5_mul2_0_1_U27 ( .A(s5_mul2_0_1_n75), .B(s5_mul2_0_1_n74), .Z(
        s5_mul2_0_1_n77) );
  XNOR2_X1 s5_mul2_0_1_U26 ( .A(s5_mul2_0_1_n73), .B(s5_mul2_0_1_n72), .ZN(
        s5_concat[14]) );
  NAND2_X1 s5_mul2_0_1_U25 ( .A1(stage4Out[6]), .A2(stage4Out[14]), .ZN(
        s5_mul2_0_1_n72) );
  XOR2_X1 s5_mul2_0_1_U24 ( .A(s5_mul2_0_1_n74), .B(s5_mul2_0_1_n71), .Z(
        s5_mul2_0_1_n73) );
  NOR2_X1 s5_mul2_0_1_U23 ( .A1(s5_mul2_0_1_n70), .A2(s5_mul2_0_1_n69), .ZN(
        s5_mul2_0_1_n74) );
  XNOR2_X1 s5_mul2_0_1_U22 ( .A(stage4Out[6]), .B(stage4Out[7]), .ZN(
        s5_mul2_0_1_n69) );
  XNOR2_X1 s5_mul2_0_1_U21 ( .A(stage4Out[14]), .B(stage4Out[15]), .ZN(
        s5_mul2_0_1_n70) );
  XNOR2_X1 s5_mul2_0_1_U20 ( .A(s5_mul2_0_1_n68), .B(s5_mul2_0_1_n67), .ZN(
        s5_concat[13]) );
  NAND2_X1 s5_mul2_0_1_U19 ( .A1(stage4Out[5]), .A2(stage4Out[13]), .ZN(
        s5_mul2_0_1_n67) );
  XOR2_X1 s5_mul2_0_1_U18 ( .A(s5_mul2_0_1_n75), .B(s5_mul2_0_1_n66), .Z(
        s5_mul2_0_1_n68) );
  XNOR2_X1 s5_mul2_0_1_U17 ( .A(s5_mul2_0_1_n65), .B(s5_mul2_0_1_n64), .ZN(
        s5_mul2_0_1_n75) );
  NAND2_X1 s5_mul2_0_1_U16 ( .A1(s5_mul2_0_1_n63), .A2(s5_mul2_0_1_n62), .ZN(
        s5_mul2_0_1_n64) );
  XNOR2_X1 s5_mul2_0_1_U15 ( .A(s5_mul2_0_1_n61), .B(s5_mul2_0_1_n60), .ZN(
        s5_mul2_0_1_n62) );
  XNOR2_X1 s5_mul2_0_1_U14 ( .A(s5_mul2_0_1_n59), .B(s5_mul2_0_1_n58), .ZN(
        s5_mul2_0_1_n63) );
  XNOR2_X1 s5_mul2_0_1_U13 ( .A(s5_mul2_0_1_n57), .B(s5_mul2_0_1_n56), .ZN(
        s5_concat[12]) );
  NAND2_X1 s5_mul2_0_1_U12 ( .A1(stage4Out[4]), .A2(stage4Out[12]), .ZN(
        s5_mul2_0_1_n56) );
  XOR2_X1 s5_mul2_0_1_U11 ( .A(s5_mul2_0_1_n66), .B(s5_mul2_0_1_n71), .Z(
        s5_mul2_0_1_n57) );
  XNOR2_X1 s5_mul2_0_1_U10 ( .A(s5_mul2_0_1_n55), .B(s5_mul2_0_1_n65), .ZN(
        s5_mul2_0_1_n71) );
  NOR2_X1 s5_mul2_0_1_U9 ( .A1(s5_mul2_0_1_n61), .A2(s5_mul2_0_1_n59), .ZN(
        s5_mul2_0_1_n65) );
  XNOR2_X1 s5_mul2_0_1_U8 ( .A(stage4Out[4]), .B(stage4Out[6]), .ZN(
        s5_mul2_0_1_n59) );
  XNOR2_X1 s5_mul2_0_1_U7 ( .A(stage4Out[12]), .B(stage4Out[14]), .ZN(
        s5_mul2_0_1_n61) );
  NAND2_X1 s5_mul2_0_1_U6 ( .A1(s5_mul2_0_1_n58), .A2(s5_mul2_0_1_n60), .ZN(
        s5_mul2_0_1_n55) );
  XOR2_X1 s5_mul2_0_1_U5 ( .A(stage4Out[13]), .B(stage4Out[15]), .Z(
        s5_mul2_0_1_n60) );
  XOR2_X1 s5_mul2_0_1_U4 ( .A(stage4Out[5]), .B(stage4Out[7]), .Z(
        s5_mul2_0_1_n58) );
  NOR2_X1 s5_mul2_0_1_U3 ( .A1(s5_mul2_0_1_n54), .A2(s5_mul2_0_1_n53), .ZN(
        s5_mul2_0_1_n66) );
  XNOR2_X1 s5_mul2_0_1_U2 ( .A(stage4Out[4]), .B(stage4Out[5]), .ZN(
        s5_mul2_0_1_n53) );
  XNOR2_X1 s5_mul2_0_1_U1 ( .A(stage4Out[12]), .B(stage4Out[13]), .ZN(
        s5_mul2_0_1_n54) );
  XNOR2_X1 s5_mul2_0_0_U29 ( .A(s5_mul2_0_0_n77), .B(s5_mul2_0_0_n76), .ZN(
        s5_concat[7]) );
  NAND2_X1 s5_mul2_0_0_U28 ( .A1(stage4Out[7]), .A2(stage4Out[3]), .ZN(
        s5_mul2_0_0_n76) );
  XOR2_X1 s5_mul2_0_0_U27 ( .A(s5_mul2_0_0_n75), .B(s5_mul2_0_0_n74), .Z(
        s5_mul2_0_0_n77) );
  XNOR2_X1 s5_mul2_0_0_U26 ( .A(s5_mul2_0_0_n73), .B(s5_mul2_0_0_n72), .ZN(
        s5_concat[6]) );
  NAND2_X1 s5_mul2_0_0_U25 ( .A1(stage4Out[6]), .A2(stage4Out[2]), .ZN(
        s5_mul2_0_0_n72) );
  XOR2_X1 s5_mul2_0_0_U24 ( .A(s5_mul2_0_0_n74), .B(s5_mul2_0_0_n71), .Z(
        s5_mul2_0_0_n73) );
  NOR2_X1 s5_mul2_0_0_U23 ( .A1(s5_mul2_0_0_n70), .A2(s5_mul2_0_0_n69), .ZN(
        s5_mul2_0_0_n74) );
  XNOR2_X1 s5_mul2_0_0_U22 ( .A(stage4Out[6]), .B(stage4Out[7]), .ZN(
        s5_mul2_0_0_n69) );
  XNOR2_X1 s5_mul2_0_0_U21 ( .A(stage4Out[2]), .B(stage4Out[3]), .ZN(
        s5_mul2_0_0_n70) );
  XNOR2_X1 s5_mul2_0_0_U20 ( .A(s5_mul2_0_0_n68), .B(s5_mul2_0_0_n67), .ZN(
        s5_concat[5]) );
  NAND2_X1 s5_mul2_0_0_U19 ( .A1(stage4Out[5]), .A2(stage4Out[1]), .ZN(
        s5_mul2_0_0_n67) );
  XOR2_X1 s5_mul2_0_0_U18 ( .A(s5_mul2_0_0_n75), .B(s5_mul2_0_0_n66), .Z(
        s5_mul2_0_0_n68) );
  XNOR2_X1 s5_mul2_0_0_U17 ( .A(s5_mul2_0_0_n65), .B(s5_mul2_0_0_n64), .ZN(
        s5_mul2_0_0_n75) );
  NAND2_X1 s5_mul2_0_0_U16 ( .A1(s5_mul2_0_0_n63), .A2(s5_mul2_0_0_n62), .ZN(
        s5_mul2_0_0_n64) );
  XNOR2_X1 s5_mul2_0_0_U15 ( .A(s5_mul2_0_0_n61), .B(s5_mul2_0_0_n60), .ZN(
        s5_mul2_0_0_n62) );
  XNOR2_X1 s5_mul2_0_0_U14 ( .A(s5_mul2_0_0_n59), .B(s5_mul2_0_0_n58), .ZN(
        s5_mul2_0_0_n63) );
  XNOR2_X1 s5_mul2_0_0_U13 ( .A(s5_mul2_0_0_n57), .B(s5_mul2_0_0_n56), .ZN(
        s5_concat[4]) );
  NAND2_X1 s5_mul2_0_0_U12 ( .A1(stage4Out[4]), .A2(stage4Out[0]), .ZN(
        s5_mul2_0_0_n56) );
  XOR2_X1 s5_mul2_0_0_U11 ( .A(s5_mul2_0_0_n66), .B(s5_mul2_0_0_n71), .Z(
        s5_mul2_0_0_n57) );
  XNOR2_X1 s5_mul2_0_0_U10 ( .A(s5_mul2_0_0_n55), .B(s5_mul2_0_0_n65), .ZN(
        s5_mul2_0_0_n71) );
  NOR2_X1 s5_mul2_0_0_U9 ( .A1(s5_mul2_0_0_n61), .A2(s5_mul2_0_0_n59), .ZN(
        s5_mul2_0_0_n65) );
  XNOR2_X1 s5_mul2_0_0_U8 ( .A(stage4Out[4]), .B(stage4Out[6]), .ZN(
        s5_mul2_0_0_n59) );
  XNOR2_X1 s5_mul2_0_0_U7 ( .A(stage4Out[0]), .B(stage4Out[2]), .ZN(
        s5_mul2_0_0_n61) );
  NAND2_X1 s5_mul2_0_0_U6 ( .A1(s5_mul2_0_0_n58), .A2(s5_mul2_0_0_n60), .ZN(
        s5_mul2_0_0_n55) );
  XOR2_X1 s5_mul2_0_0_U5 ( .A(stage4Out[1]), .B(stage4Out[3]), .Z(
        s5_mul2_0_0_n60) );
  XOR2_X1 s5_mul2_0_0_U4 ( .A(stage4Out[5]), .B(stage4Out[7]), .Z(
        s5_mul2_0_0_n58) );
  NOR2_X1 s5_mul2_0_0_U3 ( .A1(s5_mul2_0_0_n54), .A2(s5_mul2_0_0_n53), .ZN(
        s5_mul2_0_0_n66) );
  XNOR2_X1 s5_mul2_0_0_U2 ( .A(stage4Out[4]), .B(stage4Out[5]), .ZN(
        s5_mul2_0_0_n53) );
  XNOR2_X1 s5_mul2_0_0_U1 ( .A(stage4Out[0]), .B(stage4Out[1]), .ZN(
        s5_mul2_0_0_n54) );
  XOR2_X1 s5_compr_0_0_U8 ( .A(s5_regOut[7]), .B(s5_regOut[15]), .Z(
        stage5Out[7]) );
  XOR2_X1 s5_compr_0_0_U7 ( .A(s5_regOut[6]), .B(s5_regOut[14]), .Z(
        stage5Out[6]) );
  XOR2_X1 s5_compr_0_0_U6 ( .A(s5_regOut[5]), .B(s5_regOut[13]), .Z(
        stage5Out[5]) );
  XOR2_X1 s5_compr_0_0_U5 ( .A(s5_regOut[4]), .B(s5_regOut[12]), .Z(
        stage5Out[4]) );
  XOR2_X1 s5_compr_0_0_U4 ( .A(s5_regOut[3]), .B(s5_regOut[11]), .Z(
        stage5Out[3]) );
  XOR2_X1 s5_compr_0_0_U3 ( .A(s5_regOut[2]), .B(s5_regOut[10]), .Z(
        stage5Out[2]) );
  XOR2_X1 s5_compr_0_0_U2 ( .A(s5_regOut[1]), .B(s5_regOut[9]), .Z(
        stage5Out[1]) );
  XOR2_X1 s5_compr_0_0_U1 ( .A(s5_regOut[0]), .B(s5_regOut[8]), .Z(
        stage5Out[0]) );
  XOR2_X1 s5_compr_1_0_U8 ( .A(s5_regOut[23]), .B(s5_regOut[31]), .Z(
        stage5Out[15]) );
  XOR2_X1 s5_compr_1_0_U7 ( .A(s5_regOut[22]), .B(s5_regOut[30]), .Z(
        stage5Out[14]) );
  XOR2_X1 s5_compr_1_0_U6 ( .A(s5_regOut[21]), .B(s5_regOut[29]), .Z(
        stage5Out[13]) );
  XOR2_X1 s5_compr_1_0_U5 ( .A(s5_regOut[20]), .B(s5_regOut[28]), .Z(
        stage5Out[12]) );
  XOR2_X1 s5_compr_1_0_U4 ( .A(s5_regOut[19]), .B(s5_regOut[27]), .Z(
        stage5Out[11]) );
  XOR2_X1 s5_compr_1_0_U3 ( .A(s5_regOut[18]), .B(s5_regOut[26]), .Z(
        stage5Out[10]) );
  XOR2_X1 s5_compr_1_0_U2 ( .A(s5_regOut[17]), .B(s5_regOut[25]), .Z(
        stage5Out[9]) );
  XOR2_X1 s5_compr_1_0_U1 ( .A(s5_regOut[16]), .B(s5_regOut[24]), .Z(
        stage5Out[8]) );
  XOR2_X1 s6_1_U11 ( .A(stage5Out[11]), .B(stage5Out[15]), .Z(stage6Out[14])
         );
  XNOR2_X1 s6_1_U10 ( .A(stage6Out[12]), .B(s6_1_n9), .ZN(stage6Out[11]) );
  XOR2_X1 s6_1_U9 ( .A(stage6Out[15]), .B(stage5Out[15]), .Z(stage6Out[12]) );
  XNOR2_X1 s6_1_U8 ( .A(s6_1_n8), .B(stage6Out[13]), .ZN(stage6Out[10]) );
  XNOR2_X1 s6_1_U7 ( .A(stage6Out[15]), .B(stage5Out[10]), .ZN(s6_1_n8) );
  XOR2_X1 s6_1_U6 ( .A(stage5Out[14]), .B(stage5Out[8]), .Z(stage6Out[13]) );
  XOR2_X1 s6_1_U5 ( .A(stage5Out[11]), .B(stage5Out[13]), .Z(stage6Out[15]) );
  XNOR2_X1 s6_1_U4 ( .A(s6_1_n7), .B(stage5Out[9]), .ZN(stage6Out[9]) );
  XNOR2_X1 s6_1_U3 ( .A(stage5Out[13]), .B(stage5Out[12]), .ZN(s6_1_n7) );
  XNOR2_X1 s6_1_U2 ( .A(stage5Out[9]), .B(s6_1_n9), .ZN(stage6Out[8]) );
  XNOR2_X1 s6_1_U1 ( .A(stage5Out[14]), .B(stage5Out[12]), .ZN(s6_1_n9) );
  XOR2_X1 s6_0_U11 ( .A(stage5Out[3]), .B(stage5Out[7]), .Z(stage6Out[6]) );
  XNOR2_X1 s6_0_U10 ( .A(stage6Out[4]), .B(s6_0_n9), .ZN(stage6Out[3]) );
  XOR2_X1 s6_0_U9 ( .A(stage6Out[7]), .B(stage5Out[7]), .Z(stage6Out[4]) );
  XNOR2_X1 s6_0_U8 ( .A(s6_0_n8), .B(stage6Out[5]), .ZN(stage6Out[2]) );
  XNOR2_X1 s6_0_U7 ( .A(stage6Out[7]), .B(stage5Out[2]), .ZN(s6_0_n8) );
  XOR2_X1 s6_0_U6 ( .A(stage5Out[6]), .B(stage5Out[0]), .Z(stage6Out[5]) );
  XOR2_X1 s6_0_U5 ( .A(stage5Out[3]), .B(stage5Out[5]), .Z(stage6Out[7]) );
  XNOR2_X1 s6_0_U4 ( .A(s6_0_n7), .B(stage5Out[1]), .ZN(stage6Out[1]) );
  XNOR2_X1 s6_0_U3 ( .A(stage5Out[5]), .B(stage5Out[4]), .ZN(s6_0_n7) );
  XNOR2_X1 s6_0_U2 ( .A(stage5Out[1]), .B(s6_0_n9), .ZN(stage6Out[0]) );
  XNOR2_X1 s6_0_U1 ( .A(stage5Out[6]), .B(stage5Out[4]), .ZN(s6_0_n9) );
endmodule