module circuit ( clk, reset, r, input1, input2, input3, output1, output2, 
        output3, Key1, Key2, Key3, enc_dec, done );
  input [71:0] r;
  input [63:0] input1;
  input [63:0] input2;
  input [63:0] input3;
  output [63:0] output1;
  output [63:0] output2;
  output [63:0] output3;
  input [127:0] Key1;
  input [127:0] Key2;
  input [127:0] Key3;
  input clk, reset, enc_dec;
  output done;
  wire   EN, controller_n44, controller_n43, controller_n42, controller_n41,
         controller_n40, controller_n39, controller_n38, controller_n34,
         controller_n30, controller_n29, controller_n28, controller_n27,
         controller_n26, controller_n25, controller_n24, controller_n23,
         controller_n21, controller_n20, controller_n19, controller_n18,
         controller_n16, controller_n15, controller_n14, controller_n37,
         controller_n36, controller_n35, controller_n5, controller_n33,
         controller_n32, controller_n31, controller_n8, controller_n7,
         controller_N15, controller_N14, controller_N13, Midori_rounds_n2067,
         Midori_rounds_n2066, Midori_rounds_n2065, Midori_rounds_n2064,
         Midori_rounds_n2063, Midori_rounds_n2062, Midori_rounds_n2061,
         Midori_rounds_n2060, Midori_rounds_n2059, Midori_rounds_n2058,
         Midori_rounds_n2057, Midori_rounds_n2056, Midori_rounds_n2055,
         Midori_rounds_n2054, Midori_rounds_n2053, Midori_rounds_n2052,
         Midori_rounds_n2051, Midori_rounds_n2050, Midori_rounds_n2049,
         Midori_rounds_n2048, Midori_rounds_n2047, Midori_rounds_n2046,
         Midori_rounds_n2045, Midori_rounds_n2044, Midori_rounds_n2043,
         Midori_rounds_n2042, Midori_rounds_n2041, Midori_rounds_n2040,
         Midori_rounds_n2039, Midori_rounds_n2038, Midori_rounds_n2037,
         Midori_rounds_n2036, Midori_rounds_n2035, Midori_rounds_n2034,
         Midori_rounds_n2033, Midori_rounds_n2032, Midori_rounds_n2031,
         Midori_rounds_n2030, Midori_rounds_n2029, Midori_rounds_n2028,
         Midori_rounds_n2027, Midori_rounds_n2026, Midori_rounds_n2025,
         Midori_rounds_n2024, Midori_rounds_n2023, Midori_rounds_n2022,
         Midori_rounds_n2021, Midori_rounds_n2020, Midori_rounds_n2019,
         Midori_rounds_n2018, Midori_rounds_n2017, Midori_rounds_n2016,
         Midori_rounds_n2015, Midori_rounds_n2014, Midori_rounds_n2013,
         Midori_rounds_n2012, Midori_rounds_n2011, Midori_rounds_n2010,
         Midori_rounds_n2009, Midori_rounds_n2008, Midori_rounds_n2007,
         Midori_rounds_n2006, Midori_rounds_n2005, Midori_rounds_n2004,
         Midori_rounds_n2003, Midori_rounds_n2002, Midori_rounds_n2001,
         Midori_rounds_n2000, Midori_rounds_n1999, Midori_rounds_n1998,
         Midori_rounds_n1997, Midori_rounds_n1996, Midori_rounds_n1995,
         Midori_rounds_n1994, Midori_rounds_n1993, Midori_rounds_n1992,
         Midori_rounds_n1991, Midori_rounds_n1990, Midori_rounds_n1989,
         Midori_rounds_n1988, Midori_rounds_n1987, Midori_rounds_n1986,
         Midori_rounds_n1985, Midori_rounds_n1984, Midori_rounds_n1983,
         Midori_rounds_n1982, Midori_rounds_n1981, Midori_rounds_n1980,
         Midori_rounds_n1979, Midori_rounds_n1978, Midori_rounds_n1977,
         Midori_rounds_n1976, Midori_rounds_n1975, Midori_rounds_n1974,
         Midori_rounds_n1973, Midori_rounds_n1972, Midori_rounds_n1971,
         Midori_rounds_n1970, Midori_rounds_n1969, Midori_rounds_n1968,
         Midori_rounds_n1967, Midori_rounds_n1966, Midori_rounds_n1965,
         Midori_rounds_n1964, Midori_rounds_n1963, Midori_rounds_n1962,
         Midori_rounds_n1961, Midori_rounds_n1960, Midori_rounds_n1959,
         Midori_rounds_n1958, Midori_rounds_n1957, Midori_rounds_n1956,
         Midori_rounds_n1955, Midori_rounds_n1954, Midori_rounds_n1953,
         Midori_rounds_n1952, Midori_rounds_n1951, Midori_rounds_n1950,
         Midori_rounds_n1949, Midori_rounds_n1948, Midori_rounds_n1947,
         Midori_rounds_n1946, Midori_rounds_n1945, Midori_rounds_n1944,
         Midori_rounds_n1943, Midori_rounds_n1942, Midori_rounds_n1941,
         Midori_rounds_n1940, Midori_rounds_n1939, Midori_rounds_n1938,
         Midori_rounds_n1937, Midori_rounds_n1936, Midori_rounds_n1935,
         Midori_rounds_n1934, Midori_rounds_n1933, Midori_rounds_n1932,
         Midori_rounds_n1931, Midori_rounds_n1930, Midori_rounds_n1929,
         Midori_rounds_n1928, Midori_rounds_n1927, Midori_rounds_n1926,
         Midori_rounds_n1925, Midori_rounds_n1924, Midori_rounds_n1923,
         Midori_rounds_n1922, Midori_rounds_n1921, Midori_rounds_n1920,
         Midori_rounds_n1919, Midori_rounds_n1918, Midori_rounds_n1917,
         Midori_rounds_n1916, Midori_rounds_n1915, Midori_rounds_n1914,
         Midori_rounds_n1913, Midori_rounds_n1912, Midori_rounds_n1911,
         Midori_rounds_n1910, Midori_rounds_n1909, Midori_rounds_n1908,
         Midori_rounds_n1907, Midori_rounds_n1906, Midori_rounds_n1905,
         Midori_rounds_n1904, Midori_rounds_n1903, Midori_rounds_n1902,
         Midori_rounds_n1901, Midori_rounds_n1900, Midori_rounds_n1899,
         Midori_rounds_n1898, Midori_rounds_n1897, Midori_rounds_n1896,
         Midori_rounds_n1895, Midori_rounds_n1894, Midori_rounds_n1893,
         Midori_rounds_n1892, Midori_rounds_n1891, Midori_rounds_n1890,
         Midori_rounds_n1889, Midori_rounds_n1888, Midori_rounds_n1887,
         Midori_rounds_n1886, Midori_rounds_n1885, Midori_rounds_n1884,
         Midori_rounds_n1883, Midori_rounds_n1882, Midori_rounds_n1881,
         Midori_rounds_n1880, Midori_rounds_n1879, Midori_rounds_n1878,
         Midori_rounds_n1877, Midori_rounds_n1876, Midori_rounds_n1875,
         Midori_rounds_n1874, Midori_rounds_n1873, Midori_rounds_n1872,
         Midori_rounds_n1871, Midori_rounds_n1870, Midori_rounds_n1869,
         Midori_rounds_n1868, Midori_rounds_n1867, Midori_rounds_n1866,
         Midori_rounds_n1865, Midori_rounds_n1864, Midori_rounds_n1863,
         Midori_rounds_n1862, Midori_rounds_n1861, Midori_rounds_n1860,
         Midori_rounds_n1859, Midori_rounds_n1858, Midori_rounds_n1857,
         Midori_rounds_n1856, Midori_rounds_n1855, Midori_rounds_n1854,
         Midori_rounds_n1853, Midori_rounds_n1852, Midori_rounds_n1851,
         Midori_rounds_n1850, Midori_rounds_n1849, Midori_rounds_n1848,
         Midori_rounds_n1847, Midori_rounds_n1846, Midori_rounds_n1845,
         Midori_rounds_n1844, Midori_rounds_n1843, Midori_rounds_n1842,
         Midori_rounds_n1841, Midori_rounds_n1840, Midori_rounds_n1839,
         Midori_rounds_n1838, Midori_rounds_n1837, Midori_rounds_n1836,
         Midori_rounds_n1835, Midori_rounds_n1834, Midori_rounds_n1833,
         Midori_rounds_n1832, Midori_rounds_n1831, Midori_rounds_n1830,
         Midori_rounds_n1829, Midori_rounds_n1828, Midori_rounds_n1827,
         Midori_rounds_n1826, Midori_rounds_n1825, Midori_rounds_n1824,
         Midori_rounds_n1823, Midori_rounds_n1822, Midori_rounds_n1821,
         Midori_rounds_n1820, Midori_rounds_n1819, Midori_rounds_n1818,
         Midori_rounds_n1817, Midori_rounds_n1816, Midori_rounds_n1815,
         Midori_rounds_n1814, Midori_rounds_n1813, Midori_rounds_n1812,
         Midori_rounds_n1811, Midori_rounds_n1810, Midori_rounds_n1809,
         Midori_rounds_n1808, Midori_rounds_n1807, Midori_rounds_n1806,
         Midori_rounds_n1805, Midori_rounds_n1804, Midori_rounds_n1803,
         Midori_rounds_n1802, Midori_rounds_n1801, Midori_rounds_n1800,
         Midori_rounds_n1799, Midori_rounds_n1798, Midori_rounds_n1797,
         Midori_rounds_n1796, Midori_rounds_n1795, Midori_rounds_n1794,
         Midori_rounds_n1793, Midori_rounds_n1792, Midori_rounds_n1791,
         Midori_rounds_n1790, Midori_rounds_n1789, Midori_rounds_n1788,
         Midori_rounds_n1787, Midori_rounds_n1786, Midori_rounds_n1785,
         Midori_rounds_n1784, Midori_rounds_n1783, Midori_rounds_n1782,
         Midori_rounds_n1781, Midori_rounds_n1780, Midori_rounds_n1779,
         Midori_rounds_n1778, Midori_rounds_n1777, Midori_rounds_n1776,
         Midori_rounds_n1775, Midori_rounds_n1774, Midori_rounds_n1773,
         Midori_rounds_n1772, Midori_rounds_n1771, Midori_rounds_n1770,
         Midori_rounds_n1769, Midori_rounds_n1768, Midori_rounds_n1767,
         Midori_rounds_n1766, Midori_rounds_n1765, Midori_rounds_n1764,
         Midori_rounds_n1763, Midori_rounds_n1762, Midori_rounds_n1761,
         Midori_rounds_n1760, Midori_rounds_n1759, Midori_rounds_n1758,
         Midori_rounds_n1757, Midori_rounds_n1756, Midori_rounds_n1755,
         Midori_rounds_n1754, Midori_rounds_n1753, Midori_rounds_n1752,
         Midori_rounds_n1751, Midori_rounds_n1750, Midori_rounds_n1749,
         Midori_rounds_n1748, Midori_rounds_n1747, Midori_rounds_n1746,
         Midori_rounds_n1745, Midori_rounds_n1744, Midori_rounds_n1743,
         Midori_rounds_n1742, Midori_rounds_n1741, Midori_rounds_n1740,
         Midori_rounds_n1739, Midori_rounds_n1738, Midori_rounds_n1737,
         Midori_rounds_n1736, Midori_rounds_n1735, Midori_rounds_n1734,
         Midori_rounds_n1733, Midori_rounds_n1732, Midori_rounds_n1731,
         Midori_rounds_n1730, Midori_rounds_n1729, Midori_rounds_n1728,
         Midori_rounds_n1727, Midori_rounds_n1726, Midori_rounds_n1725,
         Midori_rounds_n1724, Midori_rounds_n1723, Midori_rounds_n1722,
         Midori_rounds_n1721, Midori_rounds_n1720, Midori_rounds_n1719,
         Midori_rounds_n1718, Midori_rounds_n1717, Midori_rounds_n1716,
         Midori_rounds_n1715, Midori_rounds_n1714, Midori_rounds_n1713,
         Midori_rounds_n1712, Midori_rounds_n1711, Midori_rounds_n1710,
         Midori_rounds_n1709, Midori_rounds_n1708, Midori_rounds_n1707,
         Midori_rounds_n1706, Midori_rounds_n1705, Midori_rounds_n1704,
         Midori_rounds_n1703, Midori_rounds_n1702, Midori_rounds_n1701,
         Midori_rounds_n1700, Midori_rounds_n1699, Midori_rounds_n1698,
         Midori_rounds_n1697, Midori_rounds_n1696, Midori_rounds_n1695,
         Midori_rounds_n1694, Midori_rounds_n1693, Midori_rounds_n1692,
         Midori_rounds_n1691, Midori_rounds_n1690, Midori_rounds_n1689,
         Midori_rounds_n1688, Midori_rounds_n1687, Midori_rounds_n1686,
         Midori_rounds_n1685, Midori_rounds_n1684, Midori_rounds_n1683,
         Midori_rounds_n1682, Midori_rounds_n1681, Midori_rounds_n1680,
         Midori_rounds_n1679, Midori_rounds_n1678, Midori_rounds_n1677,
         Midori_rounds_n1676, Midori_rounds_n1675, Midori_rounds_n1674,
         Midori_rounds_n1673, Midori_rounds_n1672, Midori_rounds_n1671,
         Midori_rounds_n1670, Midori_rounds_n1669, Midori_rounds_n1668,
         Midori_rounds_n1667, Midori_rounds_n1666, Midori_rounds_n1665,
         Midori_rounds_n1664, Midori_rounds_n1663, Midori_rounds_n1662,
         Midori_rounds_n1661, Midori_rounds_n1660, Midori_rounds_n1659,
         Midori_rounds_n1658, Midori_rounds_n1657, Midori_rounds_n1656,
         Midori_rounds_n1655, Midori_rounds_n1654, Midori_rounds_n1653,
         Midori_rounds_n1652, Midori_rounds_n1651, Midori_rounds_n1650,
         Midori_rounds_n1649, Midori_rounds_n1648, Midori_rounds_n1647,
         Midori_rounds_n1646, Midori_rounds_n1645, Midori_rounds_n1644,
         Midori_rounds_n1643, Midori_rounds_n1642, Midori_rounds_n1641,
         Midori_rounds_n1640, Midori_rounds_n1639, Midori_rounds_n1638,
         Midori_rounds_n1637, Midori_rounds_n1636, Midori_rounds_n1635,
         Midori_rounds_n1634, Midori_rounds_n1633, Midori_rounds_n1632,
         Midori_rounds_n1631, Midori_rounds_n1630, Midori_rounds_n1629,
         Midori_rounds_n1628, Midori_rounds_n1627, Midori_rounds_n1626,
         Midori_rounds_n1625, Midori_rounds_n1624, Midori_rounds_n1623,
         Midori_rounds_n1622, Midori_rounds_n1621, Midori_rounds_n1620,
         Midori_rounds_n1619, Midori_rounds_n1618, Midori_rounds_n1617,
         Midori_rounds_n1616, Midori_rounds_n1615, Midori_rounds_n1614,
         Midori_rounds_n1613, Midori_rounds_n1612, Midori_rounds_n1611,
         Midori_rounds_n1610, Midori_rounds_n1609, Midori_rounds_n1608,
         Midori_rounds_n1607, Midori_rounds_n1606, Midori_rounds_n1605,
         Midori_rounds_n1604, Midori_rounds_n1603, Midori_rounds_n1602,
         Midori_rounds_n1601, Midori_rounds_n1600, Midori_rounds_n1599,
         Midori_rounds_n1598, Midori_rounds_n1597, Midori_rounds_n1596,
         Midori_rounds_n1595, Midori_rounds_n1594, Midori_rounds_n1593,
         Midori_rounds_n1592, Midori_rounds_n1591, Midori_rounds_n1590,
         Midori_rounds_n1589, Midori_rounds_n1588, Midori_rounds_n1587,
         Midori_rounds_n1586, Midori_rounds_n1585, Midori_rounds_n1584,
         Midori_rounds_n1583, Midori_rounds_n1582, Midori_rounds_n1581,
         Midori_rounds_n1580, Midori_rounds_n1579, Midori_rounds_n1578,
         Midori_rounds_n1577, Midori_rounds_n1576, Midori_rounds_n1575,
         Midori_rounds_n1574, Midori_rounds_n1573, Midori_rounds_n1572,
         Midori_rounds_n1571, Midori_rounds_n1570, Midori_rounds_n1569,
         Midori_rounds_n1568, Midori_rounds_n1567, Midori_rounds_n1566,
         Midori_rounds_n1565, Midori_rounds_n1564, Midori_rounds_n1563,
         Midori_rounds_n1562, Midori_rounds_n1561, Midori_rounds_n1560,
         Midori_rounds_n1559, Midori_rounds_n1558, Midori_rounds_n1557,
         Midori_rounds_n1556, Midori_rounds_n1555, Midori_rounds_n1554,
         Midori_rounds_n1553, Midori_rounds_n1552, Midori_rounds_n1551,
         Midori_rounds_n1550, Midori_rounds_n1549, Midori_rounds_n1548,
         Midori_rounds_n1547, Midori_rounds_n1546, Midori_rounds_n1545,
         Midori_rounds_n1544, Midori_rounds_n1543, Midori_rounds_n1542,
         Midori_rounds_n1541, Midori_rounds_n1540, Midori_rounds_n1539,
         Midori_rounds_n1538, Midori_rounds_n1537, Midori_rounds_n1536,
         Midori_rounds_n1535, Midori_rounds_n1534, Midori_rounds_n1533,
         Midori_rounds_n1532, Midori_rounds_n1531, Midori_rounds_n1530,
         Midori_rounds_n1529, Midori_rounds_n1528, Midori_rounds_n1527,
         Midori_rounds_n1526, Midori_rounds_n1525, Midori_rounds_n1524,
         Midori_rounds_n1523, Midori_rounds_n1522, Midori_rounds_n1521,
         Midori_rounds_n1520, Midori_rounds_n1519, Midori_rounds_n1518,
         Midori_rounds_n1517, Midori_rounds_n1516, Midori_rounds_n1515,
         Midori_rounds_n1514, Midori_rounds_n1513, Midori_rounds_n1512,
         Midori_rounds_n1511, Midori_rounds_n1510, Midori_rounds_n1509,
         Midori_rounds_n1508, Midori_rounds_n1507, Midori_rounds_n1506,
         Midori_rounds_n1505, Midori_rounds_n1504, Midori_rounds_n1503,
         Midori_rounds_n1502, Midori_rounds_n1501, Midori_rounds_n1500,
         Midori_rounds_n1499, Midori_rounds_n1498, Midori_rounds_n1497,
         Midori_rounds_n1496, Midori_rounds_n1495, Midori_rounds_n1494,
         Midori_rounds_n1493, Midori_rounds_n1492, Midori_rounds_n1491,
         Midori_rounds_n1490, Midori_rounds_n1489, Midori_rounds_n1488,
         Midori_rounds_n1487, Midori_rounds_n1486, Midori_rounds_n1485,
         Midori_rounds_n1484, Midori_rounds_n1483, Midori_rounds_n1482,
         Midori_rounds_n1481, Midori_rounds_n1480, Midori_rounds_n1479,
         Midori_rounds_n1478, Midori_rounds_n1477, Midori_rounds_n1476,
         Midori_rounds_n1475, Midori_rounds_n1474, Midori_rounds_n1473,
         Midori_rounds_n1472, Midori_rounds_n1471, Midori_rounds_n1470,
         Midori_rounds_n1469, Midori_rounds_n1468, Midori_rounds_n1467,
         Midori_rounds_n1466, Midori_rounds_n1465, Midori_rounds_n1464,
         Midori_rounds_n1463, Midori_rounds_n1462, Midori_rounds_n1461,
         Midori_rounds_n1460, Midori_rounds_n1459, Midori_rounds_n1458,
         Midori_rounds_n1457, Midori_rounds_n1456, Midori_rounds_n1455,
         Midori_rounds_n1454, Midori_rounds_n1453, Midori_rounds_n1452,
         Midori_rounds_n1451, Midori_rounds_n1450, Midori_rounds_n1449,
         Midori_rounds_n1448, Midori_rounds_n1447, Midori_rounds_n1446,
         Midori_rounds_n1445, Midori_rounds_n1444, Midori_rounds_n1443,
         Midori_rounds_n1442, Midori_rounds_n1441, Midori_rounds_n1440,
         Midori_rounds_n1439, Midori_rounds_n1438, Midori_rounds_n1437,
         Midori_rounds_n1436, Midori_rounds_n1435, Midori_rounds_n1434,
         Midori_rounds_n1433, Midori_rounds_n1432, Midori_rounds_n1431,
         Midori_rounds_n1430, Midori_rounds_n1429, Midori_rounds_n1428,
         Midori_rounds_n1427, Midori_rounds_n1426, Midori_rounds_n1425,
         Midori_rounds_n1424, Midori_rounds_n1423, Midori_rounds_n1422,
         Midori_rounds_n1421, Midori_rounds_n1420, Midori_rounds_n1419,
         Midori_rounds_n1418, Midori_rounds_n1417, Midori_rounds_n1416,
         Midori_rounds_n1415, Midori_rounds_n1414, Midori_rounds_n1413,
         Midori_rounds_n1412, Midori_rounds_n1411, Midori_rounds_n1410,
         Midori_rounds_n1409, Midori_rounds_n1408, Midori_rounds_n1407,
         Midori_rounds_n1406, Midori_rounds_n1405, Midori_rounds_n1404,
         Midori_rounds_n1403, Midori_rounds_n1402, Midori_rounds_n1401,
         Midori_rounds_n1400, Midori_rounds_n1399, Midori_rounds_n1398,
         Midori_rounds_n1397, Midori_rounds_n1396, Midori_rounds_n1395,
         Midori_rounds_n1394, Midori_rounds_n1393, Midori_rounds_n1392,
         Midori_rounds_n1391, Midori_rounds_n1390, Midori_rounds_n1389,
         Midori_rounds_n1388, Midori_rounds_n1387, Midori_rounds_n1386,
         Midori_rounds_n1385, Midori_rounds_n1384, Midori_rounds_n1383,
         Midori_rounds_n1382, Midori_rounds_n1381, Midori_rounds_n1380,
         Midori_rounds_n1379, Midori_rounds_n1378, Midori_rounds_n1377,
         Midori_rounds_n1376, Midori_rounds_n1375, Midori_rounds_n1374,
         Midori_rounds_n1373, Midori_rounds_n1372, Midori_rounds_n1371,
         Midori_rounds_n1370, Midori_rounds_n1369, Midori_rounds_n1368,
         Midori_rounds_n1367, Midori_rounds_n1366, Midori_rounds_n1365,
         Midori_rounds_n1364, Midori_rounds_n1363, Midori_rounds_n1362,
         Midori_rounds_n1361, Midori_rounds_n1360, Midori_rounds_n1359,
         Midori_rounds_n1358, Midori_rounds_n1357, Midori_rounds_n1356,
         Midori_rounds_n1355, Midori_rounds_n1354, Midori_rounds_n1353,
         Midori_rounds_n1352, Midori_rounds_n1351, Midori_rounds_n1350,
         Midori_rounds_n1349, Midori_rounds_n1348, Midori_rounds_n1347,
         Midori_rounds_n1346, Midori_rounds_n1345, Midori_rounds_n1344,
         Midori_rounds_n1343, Midori_rounds_n1342, Midori_rounds_n1341,
         Midori_rounds_n1340, Midori_rounds_n1339, Midori_rounds_n1338,
         Midori_rounds_n1337, Midori_rounds_n1336, Midori_rounds_n1335,
         Midori_rounds_n1334, Midori_rounds_n1333, Midori_rounds_n1332,
         Midori_rounds_n1331, Midori_rounds_n1330, Midori_rounds_n1329,
         Midori_rounds_n1328, Midori_rounds_n1327, Midori_rounds_n1326,
         Midori_rounds_n1325, Midori_rounds_n1324, Midori_rounds_n1323,
         Midori_rounds_n1322, Midori_rounds_n1321, Midori_rounds_n1320,
         Midori_rounds_n1319, Midori_rounds_n1318, Midori_rounds_n1317,
         Midori_rounds_n1316, Midori_rounds_n1315, Midori_rounds_n1314,
         Midori_rounds_n1313, Midori_rounds_n1312, Midori_rounds_n1311,
         Midori_rounds_n1310, Midori_rounds_n1309, Midori_rounds_n1308,
         Midori_rounds_n1307, Midori_rounds_n1306, Midori_rounds_n1305,
         Midori_rounds_n1304, Midori_rounds_n1303, Midori_rounds_n1302,
         Midori_rounds_n1301, Midori_rounds_n1300, Midori_rounds_n1299,
         Midori_rounds_n1298, Midori_rounds_n1297, Midori_rounds_n1296,
         Midori_rounds_n1295, Midori_rounds_n1294, Midori_rounds_n1293,
         Midori_rounds_n1292, Midori_rounds_n1291, Midori_rounds_n1290,
         Midori_rounds_n1289, Midori_rounds_n1288, Midori_rounds_n1287,
         Midori_rounds_n1286, Midori_rounds_n1285, Midori_rounds_n1284,
         Midori_rounds_n1283, Midori_rounds_n1282, Midori_rounds_n1281,
         Midori_rounds_n1280, Midori_rounds_n1279, Midori_rounds_n1278,
         Midori_rounds_n1277, Midori_rounds_n1276, Midori_rounds_n1275,
         Midori_rounds_n1274, Midori_rounds_n1273, Midori_rounds_n1272,
         Midori_rounds_n1271, Midori_rounds_n1270, Midori_rounds_n1269,
         Midori_rounds_n1268, Midori_rounds_n1267, Midori_rounds_n1266,
         Midori_rounds_n1265, Midori_rounds_n1264, Midori_rounds_n1263,
         Midori_rounds_n1262, Midori_rounds_n1261, Midori_rounds_n1260,
         Midori_rounds_n1259, Midori_rounds_n1258, Midori_rounds_n1257,
         Midori_rounds_n1256, Midori_rounds_n1255, Midori_rounds_n1254,
         Midori_rounds_n1253, Midori_rounds_n1252, Midori_rounds_n1251,
         Midori_rounds_n1250, Midori_rounds_n1249, Midori_rounds_n1248,
         Midori_rounds_n1247, Midori_rounds_n1246, Midori_rounds_n1245,
         Midori_rounds_n1244, Midori_rounds_n1243, Midori_rounds_n1242,
         Midori_rounds_n1241, Midori_rounds_n979, Midori_rounds_n975,
         Midori_rounds_n971, Midori_rounds_n967, Midori_rounds_n963,
         Midori_rounds_n959, Midori_rounds_n955, Midori_rounds_n951,
         Midori_rounds_n947, Midori_rounds_n943, Midori_rounds_n939,
         Midori_rounds_n935, Midori_rounds_n931, Midori_rounds_n927,
         Midori_rounds_n923, Midori_rounds_n919, Midori_rounds_n915,
         Midori_rounds_n911, Midori_rounds_n907, Midori_rounds_n903,
         Midori_rounds_n899, Midori_rounds_n895, Midori_rounds_n891,
         Midori_rounds_n887, Midori_rounds_n883, Midori_rounds_n879,
         Midori_rounds_n875, Midori_rounds_n871, Midori_rounds_n867,
         Midori_rounds_n863, Midori_rounds_n859, Midori_rounds_n855,
         Midori_rounds_n851, Midori_rounds_n848, Midori_rounds_n845,
         Midori_rounds_n842, Midori_rounds_n839, Midori_rounds_n836,
         Midori_rounds_n833, Midori_rounds_n830, Midori_rounds_n827,
         Midori_rounds_n824, Midori_rounds_n821, Midori_rounds_n818,
         Midori_rounds_n815, Midori_rounds_n812, Midori_rounds_n809,
         Midori_rounds_n806, Midori_rounds_constant_MUX_n70,
         Midori_rounds_constant_MUX_n69, Midori_rounds_constant_MUX_n68,
         Midori_rounds_constant_MUX_n67, Midori_rounds_constant_MUX_n66,
         Midori_rounds_constant_MUX_n65, Midori_rounds_constant_MUX_n64,
         Midori_rounds_constant_MUX_n63, Midori_rounds_constant_MUX_n62,
         Midori_rounds_constant_MUX_n61, Midori_rounds_constant_MUX_n60,
         Midori_rounds_constant_MUX_n59, Midori_rounds_constant_MUX_n58,
         Midori_rounds_constant_MUX_n57, Midori_rounds_constant_MUX_n56,
         Midori_rounds_constant_MUX_n55, Midori_rounds_constant_MUX_n54,
         Midori_rounds_constant_MUX_n53, Midori_rounds_constant_MUX_n52,
         Midori_rounds_constant_MUX_n51, Midori_rounds_constant_MUX_n50,
         Midori_rounds_constant_MUX_n49, Midori_rounds_constant_MUX_n48,
         Midori_rounds_constant_MUX_n47, Midori_rounds_constant_MUX_n46,
         Midori_rounds_constant_MUX_n45, Midori_rounds_constant_MUX_n44,
         Midori_rounds_constant_MUX_n43, Midori_rounds_constant_MUX_n42,
         Midori_rounds_constant_MUX_n41, Midori_rounds_constant_MUX_n40,
         Midori_rounds_constant_MUX_n39, Midori_rounds_constant_MUX_n38,
         Midori_rounds_constant_MUX_n37, Midori_rounds_constant_MUX_n36,
         Midori_rounds_constant_MUX_n35, Midori_rounds_constant_MUX_n34,
         Midori_rounds_constant_MUX_n33, Midori_rounds_constant_MUX_n32,
         Midori_rounds_constant_MUX_n31, Midori_rounds_constant_MUX_n30,
         Midori_rounds_constant_MUX_n29, Midori_rounds_constant_MUX_n28,
         Midori_rounds_constant_MUX_n27, Midori_rounds_constant_MUX_n26,
         Midori_rounds_constant_MUX_n25, Midori_rounds_constant_MUX_n24,
         Midori_rounds_constant_MUX_n23, Midori_rounds_constant_MUX_n22,
         Midori_rounds_constant_MUX_n21, Midori_rounds_constant_MUX_n20,
         Midori_rounds_constant_MUX_n19, Midori_rounds_constant_MUX_n18,
         Midori_rounds_constant_MUX_n17, Midori_rounds_constant_MUX_n16,
         Midori_rounds_constant_MUX_n15, Midori_rounds_constant_MUX_n14,
         Midori_rounds_constant_MUX_n13, Midori_rounds_constant_MUX_n12,
         Midori_rounds_constant_MUX_n11, Midori_rounds_constant_MUX_n10,
         Midori_rounds_constant_MUX_n9,
         Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_3_,
         Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_3_,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_0__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_0__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_n16,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_3__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_3__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_n16,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_6__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_6__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_n21,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_n20,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_n19,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_n18,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_n17,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_9__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_9__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_15__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_15__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_n19,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_n18,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_n17,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_n16,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_1__Compression2_n2,
         Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_0__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_6__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_7__CF_Inst_n8,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_7__CF_Inst_n7,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_9__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_15__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_18__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_18__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_21__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_21__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_24__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_24__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_n19,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_n18,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_n17,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_n16,
         Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_3_,
         Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_3_,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_0__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_0__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_n16,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_3__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_3__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_n16,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_6__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_6__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_n21,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_n20,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_n19,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_n18,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_n17,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_9__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_9__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_15__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_15__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_n19,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_n18,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_n17,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_n16,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_1__Compression2_n2,
         Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_0__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_6__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_7__CF_Inst_n8,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_7__CF_Inst_n7,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_9__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_15__CF_Inst_n3,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_18__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_18__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_21__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_21__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_24__CF_Inst_n6,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_24__CF_Inst_n5,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_n19,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_n18,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_n17,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_n16,
         Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_3_,
         Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_3_,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_0__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_0__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_n16,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_3__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_3__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_n16,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_6__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_6__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_n21,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_n20,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_n19,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_n18,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_n17,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_9__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_9__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_15__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_15__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_n19,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_n18,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_n17,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_n16,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_1__Compression2_n2,
         Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_0__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_6__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_7__CF_Inst_n8,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_7__CF_Inst_n7,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_9__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_15__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_18__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_18__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_21__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_21__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_24__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_24__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_n19,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_n18,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_n17,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_n16,
         Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_3_,
         Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_3_,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_0__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_0__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_n16,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_3__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_3__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_n16,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_6__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_6__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_n21,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_n20,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_n19,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_n18,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_n17,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_9__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_9__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_15__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_15__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_n19,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_n18,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_n17,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_n16,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_1__Compression2_n2,
         Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_0__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_6__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_7__CF_Inst_n8,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_7__CF_Inst_n7,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_9__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_15__CF_Inst_n3,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_18__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_18__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_21__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_21__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_24__CF_Inst_n6,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_24__CF_Inst_n5,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_n19,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_n18,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_n17,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_n16,
         Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_3_,
         Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_3_,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_0__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_0__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_n16,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_3__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_3__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_n16,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_6__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_6__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_n21,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_n20,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_n19,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_n18,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_n17,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_9__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_9__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_15__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_15__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_n19,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_n18,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_n17,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_n16,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_1__Compression2_n2,
         Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_0__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_6__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_7__CF_Inst_n8,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_7__CF_Inst_n7,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_9__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_15__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_18__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_18__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_21__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_21__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_24__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_24__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_n19,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_n18,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_n17,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_n16,
         Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_3_,
         Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_3_,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_0__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_0__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_n16,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_3__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_3__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_n16,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_6__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_6__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_n21,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_n20,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_n19,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_n18,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_n17,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_9__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_9__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_15__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_15__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_n19,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_n18,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_n17,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_n16,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_1__Compression2_n2,
         Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_0__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_6__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_7__CF_Inst_n8,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_7__CF_Inst_n7,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_9__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_15__CF_Inst_n3,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_18__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_18__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_21__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_21__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_24__CF_Inst_n6,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_24__CF_Inst_n5,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_n19,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_n18,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_n17,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_n16,
         Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_3_,
         Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_3_,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_0__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_0__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_n16,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_3__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_3__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_n16,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_6__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_6__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_n21,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_n20,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_n19,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_n18,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_n17,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_9__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_9__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_15__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_15__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_n19,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_n18,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_n17,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_n16,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_1__Compression2_n2,
         Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_0__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_6__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_7__CF_Inst_n8,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_7__CF_Inst_n7,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_9__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_15__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_18__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_18__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_21__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_21__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_24__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_24__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_n19,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_n18,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_n17,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_n16,
         Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_3_,
         Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_3_,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_0__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_0__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_n16,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_3__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_3__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_n16,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_6__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_6__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_n21,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_n20,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_n19,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_n18,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_n17,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_9__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_9__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_15__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_15__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_n19,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_n18,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_n17,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_n16,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_1__Compression2_n2,
         Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_0__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_6__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_7__CF_Inst_n8,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_7__CF_Inst_n7,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_9__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_15__CF_Inst_n3,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_18__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_18__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_21__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_21__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_24__CF_Inst_n6,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_24__CF_Inst_n5,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_n19,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_n18,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_n17,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_n16,
         Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_3_,
         Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_3_,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_0__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_0__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_n16,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_3__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_3__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_n16,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_6__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_6__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_n21,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_n20,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_n19,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_n18,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_n17,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_9__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_9__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_15__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_15__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_n19,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_n18,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_n17,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_n16,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_1__Compression2_n2,
         Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_0__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_6__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_7__CF_Inst_n8,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_7__CF_Inst_n7,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_9__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_15__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_18__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_18__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_21__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_21__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_24__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_24__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_n19,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_n18,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_n17,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_n16,
         Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_3_,
         Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_3_,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_0__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_0__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_n16,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_3__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_3__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_n16,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_6__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_6__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_n21,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_n20,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_n19,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_n18,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_n17,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_9__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_9__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_15__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_15__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_n19,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_n18,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_n17,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_n16,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_1__Compression2_n2,
         Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_0__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_6__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_7__CF_Inst_n8,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_7__CF_Inst_n7,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_9__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_15__CF_Inst_n3,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_18__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_18__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_21__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_21__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_24__CF_Inst_n6,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_24__CF_Inst_n5,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_n19,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_n18,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_n17,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_n16,
         Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_3_,
         Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_3_,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_0__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_0__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_n16,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_3__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_3__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_n16,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_6__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_6__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_n21,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_n20,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_n19,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_n18,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_n17,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_9__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_9__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_15__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_15__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_n19,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_n18,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_n17,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_n16,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_1__Compression2_n2,
         Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_0__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_6__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_7__CF_Inst_n8,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_7__CF_Inst_n7,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_9__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_15__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_18__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_18__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_21__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_21__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_24__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_24__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_n19,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_n18,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_n17,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_n16,
         Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_3_,
         Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_3_,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_0__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_0__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_n16,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_3__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_3__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_n16,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_6__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_6__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_n21,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_n20,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_n19,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_n18,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_n17,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_9__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_9__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_15__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_15__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_n19,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_n18,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_n17,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_n16,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_1__Compression2_n2,
         Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_0__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_6__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_7__CF_Inst_n8,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_7__CF_Inst_n7,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_9__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_15__CF_Inst_n3,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_18__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_18__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_21__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_21__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_24__CF_Inst_n6,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_24__CF_Inst_n5,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_n19,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_n18,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_n17,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_n16,
         Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_3_,
         Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_3_,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_0__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_0__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_n16,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_3__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_3__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_n16,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_6__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_6__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_n21,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_n20,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_n19,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_n18,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_n17,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_9__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_9__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_15__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_15__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_n19,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_n18,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_n17,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_n16,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_1__Compression2_n2,
         Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_0__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_6__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_7__CF_Inst_n8,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_7__CF_Inst_n7,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_9__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_15__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_18__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_18__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_21__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_21__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_24__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_24__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_n19,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_n18,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_n17,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_n16,
         Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_3_,
         Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_3_,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_0__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_0__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_n16,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_3__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_3__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_n16,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_6__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_6__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_n21,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_n20,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_n19,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_n18,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_n17,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_9__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_9__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_15__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_15__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_n19,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_n18,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_n17,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_n16,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_1__Compression2_n2,
         Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_0__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_6__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_7__CF_Inst_n8,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_7__CF_Inst_n7,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_9__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_15__CF_Inst_n3,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_18__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_18__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_21__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_21__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_24__CF_Inst_n6,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_24__CF_Inst_n5,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_n19,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_n18,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_n17,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_n16,
         Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_3_,
         Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_3_,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_0__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_0__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_n16,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_3__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_3__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_n16,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_6__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_6__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_n21,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_n20,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_n19,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_n18,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_n17,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_9__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_9__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_15__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_15__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_n19,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_n18,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_n17,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_n16,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_1__Compression2_n2,
         Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_0__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_6__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_7__CF_Inst_n8,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_7__CF_Inst_n7,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_9__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_15__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_18__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_18__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_21__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_21__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_24__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_24__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_n19,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_n18,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_n17,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_n16,
         Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_3_,
         Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_3_,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_0__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_0__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_n16,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_3__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_3__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_n16,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_6__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_6__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_n21,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_n20,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_n19,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_n18,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_n17,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_9__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_9__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_12__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_12__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_15__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_15__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_n19,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_n18,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_n17,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_n16,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_18__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_21__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_24__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_1__Compression2_n2,
         Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_0__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_3__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_6__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_7__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_7__CF_Inst_n8,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_7__CF_Inst_n7,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_9__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_12__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_15__CF_Inst_n3,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_18__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_18__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_21__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_21__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_n14,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_n13,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_24__CF_Inst_n6,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_24__CF_Inst_n5,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_n12,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_n11,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_n10,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_n9,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_n19,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_n18,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_n17,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_n16,
         Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_n15,
         Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_0__Compression1_n3,
         Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_0__Compression2_n3,
         Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_0__Compression3_n3,
         Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_1__Compression1_n3,
         Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_1__Compression2_n3,
         Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_1__Compression3_n3,
         Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_2__Compression1_n3,
         Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_2__Compression2_n3,
         Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_2__Compression3_n3,
         Midori_rounds_mul1_MC1_n24, Midori_rounds_mul1_MC1_n23,
         Midori_rounds_mul1_MC1_n22, Midori_rounds_mul1_MC1_n21,
         Midori_rounds_mul1_MC1_n20, Midori_rounds_mul1_MC1_n19,
         Midori_rounds_mul1_MC1_n18, Midori_rounds_mul1_MC1_n17,
         Midori_rounds_mul1_MC2_n24, Midori_rounds_mul1_MC2_n23,
         Midori_rounds_mul1_MC2_n22, Midori_rounds_mul1_MC2_n21,
         Midori_rounds_mul1_MC2_n20, Midori_rounds_mul1_MC2_n19,
         Midori_rounds_mul1_MC2_n18, Midori_rounds_mul1_MC2_n17,
         Midori_rounds_mul1_MC3_n24, Midori_rounds_mul1_MC3_n23,
         Midori_rounds_mul1_MC3_n22, Midori_rounds_mul1_MC3_n21,
         Midori_rounds_mul1_MC3_n20, Midori_rounds_mul1_MC3_n19,
         Midori_rounds_mul1_MC3_n18, Midori_rounds_mul1_MC3_n17,
         Midori_rounds_mul1_MC4_n24, Midori_rounds_mul1_MC4_n23,
         Midori_rounds_mul1_MC4_n22, Midori_rounds_mul1_MC4_n21,
         Midori_rounds_mul1_MC4_n20, Midori_rounds_mul1_MC4_n19,
         Midori_rounds_mul1_MC4_n18, Midori_rounds_mul1_MC4_n17,
         Midori_rounds_mul2_MC1_n24, Midori_rounds_mul2_MC1_n23,
         Midori_rounds_mul2_MC1_n22, Midori_rounds_mul2_MC1_n21,
         Midori_rounds_mul2_MC1_n20, Midori_rounds_mul2_MC1_n19,
         Midori_rounds_mul2_MC1_n18, Midori_rounds_mul2_MC1_n17,
         Midori_rounds_mul2_MC2_n24, Midori_rounds_mul2_MC2_n23,
         Midori_rounds_mul2_MC2_n22, Midori_rounds_mul2_MC2_n21,
         Midori_rounds_mul2_MC2_n20, Midori_rounds_mul2_MC2_n19,
         Midori_rounds_mul2_MC2_n18, Midori_rounds_mul2_MC2_n17,
         Midori_rounds_mul2_MC3_n24, Midori_rounds_mul2_MC3_n23,
         Midori_rounds_mul2_MC3_n22, Midori_rounds_mul2_MC3_n21,
         Midori_rounds_mul2_MC3_n20, Midori_rounds_mul2_MC3_n19,
         Midori_rounds_mul2_MC3_n18, Midori_rounds_mul2_MC3_n17,
         Midori_rounds_mul2_MC4_n24, Midori_rounds_mul2_MC4_n23,
         Midori_rounds_mul2_MC4_n22, Midori_rounds_mul2_MC4_n21,
         Midori_rounds_mul2_MC4_n20, Midori_rounds_mul2_MC4_n19,
         Midori_rounds_mul2_MC4_n18, Midori_rounds_mul2_MC4_n17,
         Midori_rounds_mul3_MC1_n24, Midori_rounds_mul3_MC1_n23,
         Midori_rounds_mul3_MC1_n22, Midori_rounds_mul3_MC1_n21,
         Midori_rounds_mul3_MC1_n20, Midori_rounds_mul3_MC1_n19,
         Midori_rounds_mul3_MC1_n18, Midori_rounds_mul3_MC1_n17,
         Midori_rounds_mul3_MC2_n24, Midori_rounds_mul3_MC2_n23,
         Midori_rounds_mul3_MC2_n22, Midori_rounds_mul3_MC2_n21,
         Midori_rounds_mul3_MC2_n20, Midori_rounds_mul3_MC2_n19,
         Midori_rounds_mul3_MC2_n18, Midori_rounds_mul3_MC2_n17,
         Midori_rounds_mul3_MC3_n24, Midori_rounds_mul3_MC3_n23,
         Midori_rounds_mul3_MC3_n22, Midori_rounds_mul3_MC3_n21,
         Midori_rounds_mul3_MC3_n20, Midori_rounds_mul3_MC3_n19,
         Midori_rounds_mul3_MC3_n18, Midori_rounds_mul3_MC3_n17,
         Midori_rounds_mul3_MC4_n24, Midori_rounds_mul3_MC4_n23,
         Midori_rounds_mul3_MC4_n22, Midori_rounds_mul3_MC4_n21,
         Midori_rounds_mul3_MC4_n20, Midori_rounds_mul3_MC4_n19,
         Midori_rounds_mul3_MC4_n18, Midori_rounds_mul3_MC4_n17;
  wire   [63:0] wk_share1;
  wire   [63:0] wk_share2;
  wire   [63:0] wk_share3;
  wire   [3:0] round_Signal;
  wire   [63:0] Midori_add_Result_Start3;
  wire   [63:0] Midori_add_Result_Start2;
  wire   [63:0] Midori_add_Result_Start1;
  wire   [63:0] Midori_rounds_SR_Inv_Result3;
  wire   [63:0] Midori_rounds_SR_Inv_Result2;
  wire   [63:0] Midori_rounds_SR_Inv_Result1;
  wire   [63:0] Midori_rounds_mul_input3;
  wire   [63:0] Midori_rounds_mul_input2;
  wire   [63:0] Midori_rounds_mul_input1;
  wire   [63:0] Midori_rounds_SR_Result3;
  wire   [63:0] Midori_rounds_SR_Result2;
  wire   [63:0] Midori_rounds_SR_Result1;
  wire   [15:0] Midori_rounds_round_Constant;
  wire   [5:0] Midori_rounds_sub_Sub_0_rs1;
  wire   [5:0] Midori_rounds_sub_Sub_0_rs2;
  wire   [3:0] Midori_rounds_sub_Sub_0_S1_Q12_1_out3;
  wire   [3:0] Midori_rounds_sub_Sub_0_S1_Q12_1_out2;
  wire   [3:0] Midori_rounds_sub_Sub_0_S1_Q12_1_out1;
  wire   [3:0] Midori_rounds_sub_Sub_0_S1_InAff_out3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_0_S1_InAff_out3;
  wire   [3:0] Midori_rounds_sub_Sub_0_S1_InAff_out2;
  wire   [3:0] Midori_rounds_sub_Sub_0_S1_InAff_out1;
  wire   [26:0] Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_0_S2_Q12_1_out3;
  wire   [3:0] Midori_rounds_sub_Sub_0_S2_Q12_1_out2;
  wire   [3:0] Midori_rounds_sub_Sub_0_S2_Q12_1_out1;
  wire   [3:0] Midori_rounds_sub_Sub_0_S2_InAff_out3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_0_S2_InAff_out3;
  wire   [3:0] Midori_rounds_sub_Sub_0_S2_InAff_out2;
  wire   [3:0] Midori_rounds_sub_Sub_0_S2_InAff_out1;
  wire   [26:0] Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out;
  wire   [5:0] Midori_rounds_sub_Sub_1_rs1;
  wire   [5:0] Midori_rounds_sub_Sub_1_rs2;
  wire   [3:0] Midori_rounds_sub_Sub_1_S1_Q12_1_out3;
  wire   [3:0] Midori_rounds_sub_Sub_1_S1_Q12_1_out2;
  wire   [3:0] Midori_rounds_sub_Sub_1_S1_Q12_1_out1;
  wire   [3:0] Midori_rounds_sub_Sub_1_S1_InAff_out3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_1_S1_InAff_out3;
  wire   [3:0] Midori_rounds_sub_Sub_1_S1_InAff_out2;
  wire   [3:0] Midori_rounds_sub_Sub_1_S1_InAff_out1;
  wire   [26:0] Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_1_S2_Q12_1_out3;
  wire   [3:0] Midori_rounds_sub_Sub_1_S2_Q12_1_out2;
  wire   [3:0] Midori_rounds_sub_Sub_1_S2_Q12_1_out1;
  wire   [3:0] Midori_rounds_sub_Sub_1_S2_InAff_out3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_1_S2_InAff_out3;
  wire   [3:0] Midori_rounds_sub_Sub_1_S2_InAff_out2;
  wire   [3:0] Midori_rounds_sub_Sub_1_S2_InAff_out1;
  wire   [26:0] Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out;
  wire   [5:0] Midori_rounds_sub_Sub_2_rs1;
  wire   [5:0] Midori_rounds_sub_Sub_2_rs2;
  wire   [3:0] Midori_rounds_sub_Sub_2_S1_Q12_1_out3;
  wire   [3:0] Midori_rounds_sub_Sub_2_S1_Q12_1_out2;
  wire   [3:0] Midori_rounds_sub_Sub_2_S1_Q12_1_out1;
  wire   [3:0] Midori_rounds_sub_Sub_2_S1_InAff_out3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_2_S1_InAff_out3;
  wire   [3:0] Midori_rounds_sub_Sub_2_S1_InAff_out2;
  wire   [3:0] Midori_rounds_sub_Sub_2_S1_InAff_out1;
  wire   [26:0] Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_2_S2_Q12_1_out3;
  wire   [3:0] Midori_rounds_sub_Sub_2_S2_Q12_1_out2;
  wire   [3:0] Midori_rounds_sub_Sub_2_S2_Q12_1_out1;
  wire   [3:0] Midori_rounds_sub_Sub_2_S2_InAff_out3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_2_S2_InAff_out3;
  wire   [3:0] Midori_rounds_sub_Sub_2_S2_InAff_out2;
  wire   [3:0] Midori_rounds_sub_Sub_2_S2_InAff_out1;
  wire   [26:0] Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out;
  wire   [5:0] Midori_rounds_sub_Sub_3_rs1;
  wire   [5:0] Midori_rounds_sub_Sub_3_rs2;
  wire   [3:0] Midori_rounds_sub_Sub_3_S1_Q12_1_out3;
  wire   [3:0] Midori_rounds_sub_Sub_3_S1_Q12_1_out2;
  wire   [3:0] Midori_rounds_sub_Sub_3_S1_Q12_1_out1;
  wire   [3:0] Midori_rounds_sub_Sub_3_S1_InAff_out3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_3_S1_InAff_out3;
  wire   [3:0] Midori_rounds_sub_Sub_3_S1_InAff_out2;
  wire   [3:0] Midori_rounds_sub_Sub_3_S1_InAff_out1;
  wire   [26:0] Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_3_S2_Q12_1_out3;
  wire   [3:0] Midori_rounds_sub_Sub_3_S2_Q12_1_out2;
  wire   [3:0] Midori_rounds_sub_Sub_3_S2_Q12_1_out1;
  wire   [3:0] Midori_rounds_sub_Sub_3_S2_InAff_out3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_3_S2_InAff_out3;
  wire   [3:0] Midori_rounds_sub_Sub_3_S2_InAff_out2;
  wire   [3:0] Midori_rounds_sub_Sub_3_S2_InAff_out1;
  wire   [26:0] Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out;
  wire   [5:0] Midori_rounds_sub_Sub_4_rs1;
  wire   [5:0] Midori_rounds_sub_Sub_4_rs2;
  wire   [3:0] Midori_rounds_sub_Sub_4_S1_Q12_1_out3;
  wire   [3:0] Midori_rounds_sub_Sub_4_S1_Q12_1_out2;
  wire   [3:0] Midori_rounds_sub_Sub_4_S1_Q12_1_out1;
  wire   [3:0] Midori_rounds_sub_Sub_4_S1_InAff_out3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_4_S1_InAff_out3;
  wire   [3:0] Midori_rounds_sub_Sub_4_S1_InAff_out2;
  wire   [3:0] Midori_rounds_sub_Sub_4_S1_InAff_out1;
  wire   [26:0] Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_4_S2_Q12_1_out3;
  wire   [3:0] Midori_rounds_sub_Sub_4_S2_Q12_1_out2;
  wire   [3:0] Midori_rounds_sub_Sub_4_S2_Q12_1_out1;
  wire   [3:0] Midori_rounds_sub_Sub_4_S2_InAff_out3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_4_S2_InAff_out3;
  wire   [3:0] Midori_rounds_sub_Sub_4_S2_InAff_out2;
  wire   [3:0] Midori_rounds_sub_Sub_4_S2_InAff_out1;
  wire   [26:0] Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out;
  wire   [5:0] Midori_rounds_sub_Sub_5_rs1;
  wire   [5:0] Midori_rounds_sub_Sub_5_rs2;
  wire   [3:0] Midori_rounds_sub_Sub_5_S1_Q12_1_out3;
  wire   [3:0] Midori_rounds_sub_Sub_5_S1_Q12_1_out2;
  wire   [3:0] Midori_rounds_sub_Sub_5_S1_Q12_1_out1;
  wire   [3:0] Midori_rounds_sub_Sub_5_S1_InAff_out3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_5_S1_InAff_out3;
  wire   [3:0] Midori_rounds_sub_Sub_5_S1_InAff_out2;
  wire   [3:0] Midori_rounds_sub_Sub_5_S1_InAff_out1;
  wire   [26:0] Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_5_S2_Q12_1_out3;
  wire   [3:0] Midori_rounds_sub_Sub_5_S2_Q12_1_out2;
  wire   [3:0] Midori_rounds_sub_Sub_5_S2_Q12_1_out1;
  wire   [3:0] Midori_rounds_sub_Sub_5_S2_InAff_out3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_5_S2_InAff_out3;
  wire   [3:0] Midori_rounds_sub_Sub_5_S2_InAff_out2;
  wire   [3:0] Midori_rounds_sub_Sub_5_S2_InAff_out1;
  wire   [26:0] Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out;
  wire   [5:0] Midori_rounds_sub_Sub_6_rs1;
  wire   [5:0] Midori_rounds_sub_Sub_6_rs2;
  wire   [3:0] Midori_rounds_sub_Sub_6_S1_Q12_1_out3;
  wire   [3:0] Midori_rounds_sub_Sub_6_S1_Q12_1_out2;
  wire   [3:0] Midori_rounds_sub_Sub_6_S1_Q12_1_out1;
  wire   [3:0] Midori_rounds_sub_Sub_6_S1_InAff_out3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_6_S1_InAff_out3;
  wire   [3:0] Midori_rounds_sub_Sub_6_S1_InAff_out2;
  wire   [3:0] Midori_rounds_sub_Sub_6_S1_InAff_out1;
  wire   [26:0] Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_6_S2_Q12_1_out3;
  wire   [3:0] Midori_rounds_sub_Sub_6_S2_Q12_1_out2;
  wire   [3:0] Midori_rounds_sub_Sub_6_S2_Q12_1_out1;
  wire   [3:0] Midori_rounds_sub_Sub_6_S2_InAff_out3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_6_S2_InAff_out3;
  wire   [3:0] Midori_rounds_sub_Sub_6_S2_InAff_out2;
  wire   [3:0] Midori_rounds_sub_Sub_6_S2_InAff_out1;
  wire   [26:0] Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out;
  wire   [5:0] Midori_rounds_sub_Sub_7_rs1;
  wire   [5:0] Midori_rounds_sub_Sub_7_rs2;
  wire   [3:0] Midori_rounds_sub_Sub_7_S1_Q12_1_out3;
  wire   [3:0] Midori_rounds_sub_Sub_7_S1_Q12_1_out2;
  wire   [3:0] Midori_rounds_sub_Sub_7_S1_Q12_1_out1;
  wire   [3:0] Midori_rounds_sub_Sub_7_S1_InAff_out3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_7_S1_InAff_out3;
  wire   [3:0] Midori_rounds_sub_Sub_7_S1_InAff_out2;
  wire   [3:0] Midori_rounds_sub_Sub_7_S1_InAff_out1;
  wire   [26:0] Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out;
  wire   [3:0] Midori_rounds_sub_Sub_7_S2_Q12_1_out3;
  wire   [3:0] Midori_rounds_sub_Sub_7_S2_Q12_1_out2;
  wire   [3:0] Midori_rounds_sub_Sub_7_S2_Q12_1_out1;
  wire   [3:0] Midori_rounds_sub_Sub_7_S2_InAff_out3_reg;
  wire   [3:0] Midori_rounds_sub_Sub_7_S2_InAff_out3;
  wire   [3:0] Midori_rounds_sub_Sub_7_S2_InAff_out2;
  wire   [3:0] Midori_rounds_sub_Sub_7_S2_InAff_out1;
  wire   [26:0] Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out;
  wire   [26:0] Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg;
  wire   [26:0] Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out;

  XOR2_X1 KeySchadule1_U64 ( .A(Key1[73]), .B(Key1[9]), .Z(wk_share1[9]) );
  XOR2_X1 KeySchadule1_U63 ( .A(Key1[72]), .B(Key1[8]), .Z(wk_share1[8]) );
  XOR2_X1 KeySchadule1_U62 ( .A(Key1[71]), .B(Key1[7]), .Z(wk_share1[7]) );
  XOR2_X1 KeySchadule1_U61 ( .A(Key1[6]), .B(Key1[70]), .Z(wk_share1[6]) );
  XOR2_X1 KeySchadule1_U60 ( .A(Key1[127]), .B(Key1[63]), .Z(wk_share1[63]) );
  XOR2_X1 KeySchadule1_U59 ( .A(Key1[126]), .B(Key1[62]), .Z(wk_share1[62]) );
  XOR2_X1 KeySchadule1_U58 ( .A(Key1[125]), .B(Key1[61]), .Z(wk_share1[61]) );
  XOR2_X1 KeySchadule1_U57 ( .A(Key1[124]), .B(Key1[60]), .Z(wk_share1[60]) );
  XOR2_X1 KeySchadule1_U56 ( .A(Key1[5]), .B(Key1[69]), .Z(wk_share1[5]) );
  XOR2_X1 KeySchadule1_U55 ( .A(Key1[123]), .B(Key1[59]), .Z(wk_share1[59]) );
  XOR2_X1 KeySchadule1_U54 ( .A(Key1[122]), .B(Key1[58]), .Z(wk_share1[58]) );
  XOR2_X1 KeySchadule1_U53 ( .A(Key1[121]), .B(Key1[57]), .Z(wk_share1[57]) );
  XOR2_X1 KeySchadule1_U52 ( .A(Key1[120]), .B(Key1[56]), .Z(wk_share1[56]) );
  XOR2_X1 KeySchadule1_U51 ( .A(Key1[119]), .B(Key1[55]), .Z(wk_share1[55]) );
  XOR2_X1 KeySchadule1_U50 ( .A(Key1[118]), .B(Key1[54]), .Z(wk_share1[54]) );
  XOR2_X1 KeySchadule1_U49 ( .A(Key1[117]), .B(Key1[53]), .Z(wk_share1[53]) );
  XOR2_X1 KeySchadule1_U48 ( .A(Key1[116]), .B(Key1[52]), .Z(wk_share1[52]) );
  XOR2_X1 KeySchadule1_U47 ( .A(Key1[115]), .B(Key1[51]), .Z(wk_share1[51]) );
  XOR2_X1 KeySchadule1_U46 ( .A(Key1[114]), .B(Key1[50]), .Z(wk_share1[50]) );
  XOR2_X1 KeySchadule1_U45 ( .A(Key1[4]), .B(Key1[68]), .Z(wk_share1[4]) );
  XOR2_X1 KeySchadule1_U44 ( .A(Key1[113]), .B(Key1[49]), .Z(wk_share1[49]) );
  XOR2_X1 KeySchadule1_U43 ( .A(Key1[112]), .B(Key1[48]), .Z(wk_share1[48]) );
  XOR2_X1 KeySchadule1_U42 ( .A(Key1[111]), .B(Key1[47]), .Z(wk_share1[47]) );
  XOR2_X1 KeySchadule1_U41 ( .A(Key1[110]), .B(Key1[46]), .Z(wk_share1[46]) );
  XOR2_X1 KeySchadule1_U40 ( .A(Key1[109]), .B(Key1[45]), .Z(wk_share1[45]) );
  XOR2_X1 KeySchadule1_U39 ( .A(Key1[108]), .B(Key1[44]), .Z(wk_share1[44]) );
  XOR2_X1 KeySchadule1_U38 ( .A(Key1[107]), .B(Key1[43]), .Z(wk_share1[43]) );
  XOR2_X1 KeySchadule1_U37 ( .A(Key1[106]), .B(Key1[42]), .Z(wk_share1[42]) );
  XOR2_X1 KeySchadule1_U36 ( .A(Key1[105]), .B(Key1[41]), .Z(wk_share1[41]) );
  XOR2_X1 KeySchadule1_U35 ( .A(Key1[104]), .B(Key1[40]), .Z(wk_share1[40]) );
  XOR2_X1 KeySchadule1_U34 ( .A(Key1[3]), .B(Key1[67]), .Z(wk_share1[3]) );
  XOR2_X1 KeySchadule1_U33 ( .A(Key1[103]), .B(Key1[39]), .Z(wk_share1[39]) );
  XOR2_X1 KeySchadule1_U32 ( .A(Key1[102]), .B(Key1[38]), .Z(wk_share1[38]) );
  XOR2_X1 KeySchadule1_U31 ( .A(Key1[101]), .B(Key1[37]), .Z(wk_share1[37]) );
  XOR2_X1 KeySchadule1_U30 ( .A(Key1[100]), .B(Key1[36]), .Z(wk_share1[36]) );
  XOR2_X1 KeySchadule1_U29 ( .A(Key1[35]), .B(Key1[99]), .Z(wk_share1[35]) );
  XOR2_X1 KeySchadule1_U28 ( .A(Key1[34]), .B(Key1[98]), .Z(wk_share1[34]) );
  XOR2_X1 KeySchadule1_U27 ( .A(Key1[33]), .B(Key1[97]), .Z(wk_share1[33]) );
  XOR2_X1 KeySchadule1_U26 ( .A(Key1[32]), .B(Key1[96]), .Z(wk_share1[32]) );
  XOR2_X1 KeySchadule1_U25 ( .A(Key1[31]), .B(Key1[95]), .Z(wk_share1[31]) );
  XOR2_X1 KeySchadule1_U24 ( .A(Key1[30]), .B(Key1[94]), .Z(wk_share1[30]) );
  XOR2_X1 KeySchadule1_U23 ( .A(Key1[2]), .B(Key1[66]), .Z(wk_share1[2]) );
  XOR2_X1 KeySchadule1_U22 ( .A(Key1[29]), .B(Key1[93]), .Z(wk_share1[29]) );
  XOR2_X1 KeySchadule1_U21 ( .A(Key1[28]), .B(Key1[92]), .Z(wk_share1[28]) );
  XOR2_X1 KeySchadule1_U20 ( .A(Key1[27]), .B(Key1[91]), .Z(wk_share1[27]) );
  XOR2_X1 KeySchadule1_U19 ( .A(Key1[26]), .B(Key1[90]), .Z(wk_share1[26]) );
  XOR2_X1 KeySchadule1_U18 ( .A(Key1[25]), .B(Key1[89]), .Z(wk_share1[25]) );
  XOR2_X1 KeySchadule1_U17 ( .A(Key1[24]), .B(Key1[88]), .Z(wk_share1[24]) );
  XOR2_X1 KeySchadule1_U16 ( .A(Key1[23]), .B(Key1[87]), .Z(wk_share1[23]) );
  XOR2_X1 KeySchadule1_U15 ( .A(Key1[22]), .B(Key1[86]), .Z(wk_share1[22]) );
  XOR2_X1 KeySchadule1_U14 ( .A(Key1[21]), .B(Key1[85]), .Z(wk_share1[21]) );
  XOR2_X1 KeySchadule1_U13 ( .A(Key1[20]), .B(Key1[84]), .Z(wk_share1[20]) );
  XOR2_X1 KeySchadule1_U12 ( .A(Key1[1]), .B(Key1[65]), .Z(wk_share1[1]) );
  XOR2_X1 KeySchadule1_U11 ( .A(Key1[19]), .B(Key1[83]), .Z(wk_share1[19]) );
  XOR2_X1 KeySchadule1_U10 ( .A(Key1[18]), .B(Key1[82]), .Z(wk_share1[18]) );
  XOR2_X1 KeySchadule1_U9 ( .A(Key1[17]), .B(Key1[81]), .Z(wk_share1[17]) );
  XOR2_X1 KeySchadule1_U8 ( .A(Key1[16]), .B(Key1[80]), .Z(wk_share1[16]) );
  XOR2_X1 KeySchadule1_U7 ( .A(Key1[15]), .B(Key1[79]), .Z(wk_share1[15]) );
  XOR2_X1 KeySchadule1_U6 ( .A(Key1[14]), .B(Key1[78]), .Z(wk_share1[14]) );
  XOR2_X1 KeySchadule1_U5 ( .A(Key1[13]), .B(Key1[77]), .Z(wk_share1[13]) );
  XOR2_X1 KeySchadule1_U4 ( .A(Key1[12]), .B(Key1[76]), .Z(wk_share1[12]) );
  XOR2_X1 KeySchadule1_U3 ( .A(Key1[11]), .B(Key1[75]), .Z(wk_share1[11]) );
  XOR2_X1 KeySchadule1_U2 ( .A(Key1[10]), .B(Key1[74]), .Z(wk_share1[10]) );
  XOR2_X1 KeySchadule1_U1 ( .A(Key1[0]), .B(Key1[64]), .Z(wk_share1[0]) );
  XOR2_X1 KeySchadule2_U64 ( .A(Key2[73]), .B(Key2[9]), .Z(wk_share2[9]) );
  XOR2_X1 KeySchadule2_U63 ( .A(Key2[72]), .B(Key2[8]), .Z(wk_share2[8]) );
  XOR2_X1 KeySchadule2_U62 ( .A(Key2[71]), .B(Key2[7]), .Z(wk_share2[7]) );
  XOR2_X1 KeySchadule2_U61 ( .A(Key2[6]), .B(Key2[70]), .Z(wk_share2[6]) );
  XOR2_X1 KeySchadule2_U60 ( .A(Key2[127]), .B(Key2[63]), .Z(wk_share2[63]) );
  XOR2_X1 KeySchadule2_U59 ( .A(Key2[126]), .B(Key2[62]), .Z(wk_share2[62]) );
  XOR2_X1 KeySchadule2_U58 ( .A(Key2[125]), .B(Key2[61]), .Z(wk_share2[61]) );
  XOR2_X1 KeySchadule2_U57 ( .A(Key2[124]), .B(Key2[60]), .Z(wk_share2[60]) );
  XOR2_X1 KeySchadule2_U56 ( .A(Key2[5]), .B(Key2[69]), .Z(wk_share2[5]) );
  XOR2_X1 KeySchadule2_U55 ( .A(Key2[123]), .B(Key2[59]), .Z(wk_share2[59]) );
  XOR2_X1 KeySchadule2_U54 ( .A(Key2[122]), .B(Key2[58]), .Z(wk_share2[58]) );
  XOR2_X1 KeySchadule2_U53 ( .A(Key2[121]), .B(Key2[57]), .Z(wk_share2[57]) );
  XOR2_X1 KeySchadule2_U52 ( .A(Key2[120]), .B(Key2[56]), .Z(wk_share2[56]) );
  XOR2_X1 KeySchadule2_U51 ( .A(Key2[119]), .B(Key2[55]), .Z(wk_share2[55]) );
  XOR2_X1 KeySchadule2_U50 ( .A(Key2[118]), .B(Key2[54]), .Z(wk_share2[54]) );
  XOR2_X1 KeySchadule2_U49 ( .A(Key2[117]), .B(Key2[53]), .Z(wk_share2[53]) );
  XOR2_X1 KeySchadule2_U48 ( .A(Key2[116]), .B(Key2[52]), .Z(wk_share2[52]) );
  XOR2_X1 KeySchadule2_U47 ( .A(Key2[115]), .B(Key2[51]), .Z(wk_share2[51]) );
  XOR2_X1 KeySchadule2_U46 ( .A(Key2[114]), .B(Key2[50]), .Z(wk_share2[50]) );
  XOR2_X1 KeySchadule2_U45 ( .A(Key2[4]), .B(Key2[68]), .Z(wk_share2[4]) );
  XOR2_X1 KeySchadule2_U44 ( .A(Key2[113]), .B(Key2[49]), .Z(wk_share2[49]) );
  XOR2_X1 KeySchadule2_U43 ( .A(Key2[112]), .B(Key2[48]), .Z(wk_share2[48]) );
  XOR2_X1 KeySchadule2_U42 ( .A(Key2[111]), .B(Key2[47]), .Z(wk_share2[47]) );
  XOR2_X1 KeySchadule2_U41 ( .A(Key2[110]), .B(Key2[46]), .Z(wk_share2[46]) );
  XOR2_X1 KeySchadule2_U40 ( .A(Key2[109]), .B(Key2[45]), .Z(wk_share2[45]) );
  XOR2_X1 KeySchadule2_U39 ( .A(Key2[108]), .B(Key2[44]), .Z(wk_share2[44]) );
  XOR2_X1 KeySchadule2_U38 ( .A(Key2[107]), .B(Key2[43]), .Z(wk_share2[43]) );
  XOR2_X1 KeySchadule2_U37 ( .A(Key2[106]), .B(Key2[42]), .Z(wk_share2[42]) );
  XOR2_X1 KeySchadule2_U36 ( .A(Key2[105]), .B(Key2[41]), .Z(wk_share2[41]) );
  XOR2_X1 KeySchadule2_U35 ( .A(Key2[104]), .B(Key2[40]), .Z(wk_share2[40]) );
  XOR2_X1 KeySchadule2_U34 ( .A(Key2[3]), .B(Key2[67]), .Z(wk_share2[3]) );
  XOR2_X1 KeySchadule2_U33 ( .A(Key2[103]), .B(Key2[39]), .Z(wk_share2[39]) );
  XOR2_X1 KeySchadule2_U32 ( .A(Key2[102]), .B(Key2[38]), .Z(wk_share2[38]) );
  XOR2_X1 KeySchadule2_U31 ( .A(Key2[101]), .B(Key2[37]), .Z(wk_share2[37]) );
  XOR2_X1 KeySchadule2_U30 ( .A(Key2[100]), .B(Key2[36]), .Z(wk_share2[36]) );
  XOR2_X1 KeySchadule2_U29 ( .A(Key2[35]), .B(Key2[99]), .Z(wk_share2[35]) );
  XOR2_X1 KeySchadule2_U28 ( .A(Key2[34]), .B(Key2[98]), .Z(wk_share2[34]) );
  XOR2_X1 KeySchadule2_U27 ( .A(Key2[33]), .B(Key2[97]), .Z(wk_share2[33]) );
  XOR2_X1 KeySchadule2_U26 ( .A(Key2[32]), .B(Key2[96]), .Z(wk_share2[32]) );
  XOR2_X1 KeySchadule2_U25 ( .A(Key2[31]), .B(Key2[95]), .Z(wk_share2[31]) );
  XOR2_X1 KeySchadule2_U24 ( .A(Key2[30]), .B(Key2[94]), .Z(wk_share2[30]) );
  XOR2_X1 KeySchadule2_U23 ( .A(Key2[2]), .B(Key2[66]), .Z(wk_share2[2]) );
  XOR2_X1 KeySchadule2_U22 ( .A(Key2[29]), .B(Key2[93]), .Z(wk_share2[29]) );
  XOR2_X1 KeySchadule2_U21 ( .A(Key2[28]), .B(Key2[92]), .Z(wk_share2[28]) );
  XOR2_X1 KeySchadule2_U20 ( .A(Key2[27]), .B(Key2[91]), .Z(wk_share2[27]) );
  XOR2_X1 KeySchadule2_U19 ( .A(Key2[26]), .B(Key2[90]), .Z(wk_share2[26]) );
  XOR2_X1 KeySchadule2_U18 ( .A(Key2[25]), .B(Key2[89]), .Z(wk_share2[25]) );
  XOR2_X1 KeySchadule2_U17 ( .A(Key2[24]), .B(Key2[88]), .Z(wk_share2[24]) );
  XOR2_X1 KeySchadule2_U16 ( .A(Key2[23]), .B(Key2[87]), .Z(wk_share2[23]) );
  XOR2_X1 KeySchadule2_U15 ( .A(Key2[22]), .B(Key2[86]), .Z(wk_share2[22]) );
  XOR2_X1 KeySchadule2_U14 ( .A(Key2[21]), .B(Key2[85]), .Z(wk_share2[21]) );
  XOR2_X1 KeySchadule2_U13 ( .A(Key2[20]), .B(Key2[84]), .Z(wk_share2[20]) );
  XOR2_X1 KeySchadule2_U12 ( .A(Key2[1]), .B(Key2[65]), .Z(wk_share2[1]) );
  XOR2_X1 KeySchadule2_U11 ( .A(Key2[19]), .B(Key2[83]), .Z(wk_share2[19]) );
  XOR2_X1 KeySchadule2_U10 ( .A(Key2[18]), .B(Key2[82]), .Z(wk_share2[18]) );
  XOR2_X1 KeySchadule2_U9 ( .A(Key2[17]), .B(Key2[81]), .Z(wk_share2[17]) );
  XOR2_X1 KeySchadule2_U8 ( .A(Key2[16]), .B(Key2[80]), .Z(wk_share2[16]) );
  XOR2_X1 KeySchadule2_U7 ( .A(Key2[15]), .B(Key2[79]), .Z(wk_share2[15]) );
  XOR2_X1 KeySchadule2_U6 ( .A(Key2[14]), .B(Key2[78]), .Z(wk_share2[14]) );
  XOR2_X1 KeySchadule2_U5 ( .A(Key2[13]), .B(Key2[77]), .Z(wk_share2[13]) );
  XOR2_X1 KeySchadule2_U4 ( .A(Key2[12]), .B(Key2[76]), .Z(wk_share2[12]) );
  XOR2_X1 KeySchadule2_U3 ( .A(Key2[11]), .B(Key2[75]), .Z(wk_share2[11]) );
  XOR2_X1 KeySchadule2_U2 ( .A(Key2[10]), .B(Key2[74]), .Z(wk_share2[10]) );
  XOR2_X1 KeySchadule2_U1 ( .A(Key2[0]), .B(Key2[64]), .Z(wk_share2[0]) );
  XOR2_X1 KeySchadule3_U64 ( .A(Key3[73]), .B(Key3[9]), .Z(wk_share3[9]) );
  XOR2_X1 KeySchadule3_U63 ( .A(Key3[72]), .B(Key3[8]), .Z(wk_share3[8]) );
  XOR2_X1 KeySchadule3_U62 ( .A(Key3[71]), .B(Key3[7]), .Z(wk_share3[7]) );
  XOR2_X1 KeySchadule3_U61 ( .A(Key3[6]), .B(Key3[70]), .Z(wk_share3[6]) );
  XOR2_X1 KeySchadule3_U60 ( .A(Key3[127]), .B(Key3[63]), .Z(wk_share3[63]) );
  XOR2_X1 KeySchadule3_U59 ( .A(Key3[126]), .B(Key3[62]), .Z(wk_share3[62]) );
  XOR2_X1 KeySchadule3_U58 ( .A(Key3[125]), .B(Key3[61]), .Z(wk_share3[61]) );
  XOR2_X1 KeySchadule3_U57 ( .A(Key3[124]), .B(Key3[60]), .Z(wk_share3[60]) );
  XOR2_X1 KeySchadule3_U56 ( .A(Key3[5]), .B(Key3[69]), .Z(wk_share3[5]) );
  XOR2_X1 KeySchadule3_U55 ( .A(Key3[123]), .B(Key3[59]), .Z(wk_share3[59]) );
  XOR2_X1 KeySchadule3_U54 ( .A(Key3[122]), .B(Key3[58]), .Z(wk_share3[58]) );
  XOR2_X1 KeySchadule3_U53 ( .A(Key3[121]), .B(Key3[57]), .Z(wk_share3[57]) );
  XOR2_X1 KeySchadule3_U52 ( .A(Key3[120]), .B(Key3[56]), .Z(wk_share3[56]) );
  XOR2_X1 KeySchadule3_U51 ( .A(Key3[119]), .B(Key3[55]), .Z(wk_share3[55]) );
  XOR2_X1 KeySchadule3_U50 ( .A(Key3[118]), .B(Key3[54]), .Z(wk_share3[54]) );
  XOR2_X1 KeySchadule3_U49 ( .A(Key3[117]), .B(Key3[53]), .Z(wk_share3[53]) );
  XOR2_X1 KeySchadule3_U48 ( .A(Key3[116]), .B(Key3[52]), .Z(wk_share3[52]) );
  XOR2_X1 KeySchadule3_U47 ( .A(Key3[115]), .B(Key3[51]), .Z(wk_share3[51]) );
  XOR2_X1 KeySchadule3_U46 ( .A(Key3[114]), .B(Key3[50]), .Z(wk_share3[50]) );
  XOR2_X1 KeySchadule3_U45 ( .A(Key3[4]), .B(Key3[68]), .Z(wk_share3[4]) );
  XOR2_X1 KeySchadule3_U44 ( .A(Key3[113]), .B(Key3[49]), .Z(wk_share3[49]) );
  XOR2_X1 KeySchadule3_U43 ( .A(Key3[112]), .B(Key3[48]), .Z(wk_share3[48]) );
  XOR2_X1 KeySchadule3_U42 ( .A(Key3[111]), .B(Key3[47]), .Z(wk_share3[47]) );
  XOR2_X1 KeySchadule3_U41 ( .A(Key3[110]), .B(Key3[46]), .Z(wk_share3[46]) );
  XOR2_X1 KeySchadule3_U40 ( .A(Key3[109]), .B(Key3[45]), .Z(wk_share3[45]) );
  XOR2_X1 KeySchadule3_U39 ( .A(Key3[108]), .B(Key3[44]), .Z(wk_share3[44]) );
  XOR2_X1 KeySchadule3_U38 ( .A(Key3[107]), .B(Key3[43]), .Z(wk_share3[43]) );
  XOR2_X1 KeySchadule3_U37 ( .A(Key3[106]), .B(Key3[42]), .Z(wk_share3[42]) );
  XOR2_X1 KeySchadule3_U36 ( .A(Key3[105]), .B(Key3[41]), .Z(wk_share3[41]) );
  XOR2_X1 KeySchadule3_U35 ( .A(Key3[104]), .B(Key3[40]), .Z(wk_share3[40]) );
  XOR2_X1 KeySchadule3_U34 ( .A(Key3[3]), .B(Key3[67]), .Z(wk_share3[3]) );
  XOR2_X1 KeySchadule3_U33 ( .A(Key3[103]), .B(Key3[39]), .Z(wk_share3[39]) );
  XOR2_X1 KeySchadule3_U32 ( .A(Key3[102]), .B(Key3[38]), .Z(wk_share3[38]) );
  XOR2_X1 KeySchadule3_U31 ( .A(Key3[101]), .B(Key3[37]), .Z(wk_share3[37]) );
  XOR2_X1 KeySchadule3_U30 ( .A(Key3[100]), .B(Key3[36]), .Z(wk_share3[36]) );
  XOR2_X1 KeySchadule3_U29 ( .A(Key3[35]), .B(Key3[99]), .Z(wk_share3[35]) );
  XOR2_X1 KeySchadule3_U28 ( .A(Key3[34]), .B(Key3[98]), .Z(wk_share3[34]) );
  XOR2_X1 KeySchadule3_U27 ( .A(Key3[33]), .B(Key3[97]), .Z(wk_share3[33]) );
  XOR2_X1 KeySchadule3_U26 ( .A(Key3[32]), .B(Key3[96]), .Z(wk_share3[32]) );
  XOR2_X1 KeySchadule3_U25 ( .A(Key3[31]), .B(Key3[95]), .Z(wk_share3[31]) );
  XOR2_X1 KeySchadule3_U24 ( .A(Key3[30]), .B(Key3[94]), .Z(wk_share3[30]) );
  XOR2_X1 KeySchadule3_U23 ( .A(Key3[2]), .B(Key3[66]), .Z(wk_share3[2]) );
  XOR2_X1 KeySchadule3_U22 ( .A(Key3[29]), .B(Key3[93]), .Z(wk_share3[29]) );
  XOR2_X1 KeySchadule3_U21 ( .A(Key3[28]), .B(Key3[92]), .Z(wk_share3[28]) );
  XOR2_X1 KeySchadule3_U20 ( .A(Key3[27]), .B(Key3[91]), .Z(wk_share3[27]) );
  XOR2_X1 KeySchadule3_U19 ( .A(Key3[26]), .B(Key3[90]), .Z(wk_share3[26]) );
  XOR2_X1 KeySchadule3_U18 ( .A(Key3[25]), .B(Key3[89]), .Z(wk_share3[25]) );
  XOR2_X1 KeySchadule3_U17 ( .A(Key3[24]), .B(Key3[88]), .Z(wk_share3[24]) );
  XOR2_X1 KeySchadule3_U16 ( .A(Key3[23]), .B(Key3[87]), .Z(wk_share3[23]) );
  XOR2_X1 KeySchadule3_U15 ( .A(Key3[22]), .B(Key3[86]), .Z(wk_share3[22]) );
  XOR2_X1 KeySchadule3_U14 ( .A(Key3[21]), .B(Key3[85]), .Z(wk_share3[21]) );
  XOR2_X1 KeySchadule3_U13 ( .A(Key3[20]), .B(Key3[84]), .Z(wk_share3[20]) );
  XOR2_X1 KeySchadule3_U12 ( .A(Key3[1]), .B(Key3[65]), .Z(wk_share3[1]) );
  XOR2_X1 KeySchadule3_U11 ( .A(Key3[19]), .B(Key3[83]), .Z(wk_share3[19]) );
  XOR2_X1 KeySchadule3_U10 ( .A(Key3[18]), .B(Key3[82]), .Z(wk_share3[18]) );
  XOR2_X1 KeySchadule3_U9 ( .A(Key3[17]), .B(Key3[81]), .Z(wk_share3[17]) );
  XOR2_X1 KeySchadule3_U8 ( .A(Key3[16]), .B(Key3[80]), .Z(wk_share3[16]) );
  XOR2_X1 KeySchadule3_U7 ( .A(Key3[15]), .B(Key3[79]), .Z(wk_share3[15]) );
  XOR2_X1 KeySchadule3_U6 ( .A(Key3[14]), .B(Key3[78]), .Z(wk_share3[14]) );
  XOR2_X1 KeySchadule3_U5 ( .A(Key3[13]), .B(Key3[77]), .Z(wk_share3[13]) );
  XOR2_X1 KeySchadule3_U4 ( .A(Key3[12]), .B(Key3[76]), .Z(wk_share3[12]) );
  XOR2_X1 KeySchadule3_U3 ( .A(Key3[11]), .B(Key3[75]), .Z(wk_share3[11]) );
  XOR2_X1 KeySchadule3_U2 ( .A(Key3[10]), .B(Key3[74]), .Z(wk_share3[10]) );
  XOR2_X1 KeySchadule3_U1 ( .A(Key3[0]), .B(Key3[64]), .Z(wk_share3[0]) );
  AOI22_X1 controller_U32 ( .A1(round_Signal[0]), .A2(controller_n44), .B1(
        controller_n43), .B2(controller_n18), .ZN(controller_n33) );
  INV_X1 controller_U31 ( .A(controller_n42), .ZN(controller_n32) );
  AOI22_X1 controller_U30 ( .A1(round_Signal[2]), .A2(controller_n41), .B1(
        controller_n40), .B2(controller_n39), .ZN(controller_n42) );
  NOR2_X1 controller_U29 ( .A1(controller_n18), .A2(controller_n20), .ZN(
        controller_n39) );
  AOI22_X1 controller_U28 ( .A1(round_Signal[1]), .A2(controller_n38), .B1(
        controller_n34), .B2(controller_n20), .ZN(controller_n5) );
  OAI22_X1 controller_U27 ( .A1(controller_n36), .A2(controller_n30), .B1(
        reset), .B2(controller_n29), .ZN(controller_n37) );
  OAI221_X1 controller_U26 ( .B1(controller_n7), .B2(controller_n36), .C1(
        controller_n7), .C2(controller_n28), .A(controller_n27), .ZN(
        controller_n29) );
  OAI21_X1 controller_U25 ( .B1(round_Signal[1]), .B2(controller_n43), .A(
        controller_n38), .ZN(controller_n41) );
  NAND2_X1 controller_U24 ( .A1(controller_n23), .A2(controller_n34), .ZN(
        controller_n38) );
  OR2_X1 controller_U23 ( .A1(controller_n43), .A2(controller_n18), .ZN(
        controller_n34) );
  NOR2_X1 controller_U22 ( .A1(round_Signal[2]), .A2(controller_n43), .ZN(
        controller_n40) );
  NAND2_X1 controller_U21 ( .A1(controller_n25), .A2(controller_n23), .ZN(
        controller_n43) );
  AOI21_X1 controller_U20 ( .B1(controller_n8), .B2(controller_n23), .A(
        controller_N13), .ZN(controller_n30) );
  AOI211_X1 controller_U19 ( .C1(controller_n35), .C2(controller_n8), .A(
        controller_n28), .B(controller_n44), .ZN(controller_N14) );
  NOR2_X1 controller_U18 ( .A1(controller_n21), .A2(controller_n44), .ZN(
        controller_N13) );
  NOR3_X1 controller_U17 ( .A1(controller_n8), .A2(controller_n27), .A3(
        controller_n21), .ZN(controller_n25) );
  NAND3_X1 controller_U16 ( .A1(controller_n24), .A2(controller_n28), .A3(done), .ZN(EN) );
  NOR2_X1 controller_U15 ( .A1(controller_n8), .A2(controller_n35), .ZN(
        controller_n28) );
  INV_X1 controller_U14 ( .A(controller_n27), .ZN(controller_n24) );
  NAND2_X1 controller_U13 ( .A1(controller_n36), .A2(controller_n7), .ZN(
        controller_n27) );
  NOR2_X1 controller_U12 ( .A1(controller_n19), .A2(controller_n26), .ZN(done)
         );
  NAND3_X1 controller_U11 ( .A1(round_Signal[2]), .A2(round_Signal[0]), .A3(
        round_Signal[1]), .ZN(controller_n26) );
  INV_X1 controller_U10 ( .A(reset), .ZN(controller_n23) );
  OR2_X1 controller_U9 ( .A1(reset), .A2(controller_n25), .ZN(controller_n44)
         );
  INV_X1 controller_U7 ( .A(controller_n19), .ZN(controller_n16) );
  NOR2_X1 controller_U6 ( .A1(controller_n41), .A2(controller_n40), .ZN(
        controller_n15) );
  OAI22_X1 controller_U5 ( .A1(controller_n44), .A2(controller_n14), .B1(
        controller_n30), .B2(controller_n7), .ZN(controller_N15) );
  NAND2_X1 controller_U4 ( .A1(controller_n7), .A2(controller_n28), .ZN(
        controller_n14) );
  OAI33_X1 controller_U3 ( .A1(1'b0), .A2(controller_n19), .A3(controller_n15), 
        .B1(controller_n16), .B2(controller_n43), .B3(controller_n26), .ZN(
        controller_n31) );
  DFF_X1 controller_PerRoundCounter_reg_2_ ( .D(controller_N15), .CK(clk), 
        .Q(), .QN(controller_n7) );
  DFF_X1 controller_PerRoundCounter_reg_3_ ( .D(controller_n37), .CK(clk), 
        .Q(), .QN(controller_n36) );
  DFF_X1 controller_RoundCounter_reg_0_ ( .D(controller_n33), .CK(clk), .Q(
        round_Signal[0]), .QN(controller_n18) );
  DFF_X1 controller_PerRoundCounter_reg_1_ ( .D(controller_N14), .CK(clk), 
        .Q(), .QN(controller_n8) );
  DFF_X1 controller_RoundCounter_reg_3_ ( .D(controller_n31), .CK(clk), .Q(
        round_Signal[3]), .QN(controller_n19) );
  DFF_X1 controller_RoundCounter_reg_2_ ( .D(controller_n32), .CK(clk), .Q(
        round_Signal[2]), .QN() );
  DFF_X1 controller_RoundCounter_reg_1_ ( .D(controller_n5), .CK(clk), .Q(
        round_Signal[1]), .QN(controller_n20) );
  DFF_X1 controller_PerRoundCounter_reg_0_ ( .D(controller_N13), .CK(clk), .Q(
        controller_n21), .QN(controller_n35) );
  XOR2_X1 Midori_U384 ( .A(wk_share3[9]), .B(Midori_rounds_SR_Result3[9]), .Z(
        output3[9]) );
  XOR2_X1 Midori_U383 ( .A(wk_share3[8]), .B(Midori_rounds_SR_Result3[8]), .Z(
        output3[8]) );
  XOR2_X1 Midori_U382 ( .A(wk_share3[7]), .B(Midori_rounds_SR_Result3[47]), 
        .Z(output3[7]) );
  XOR2_X1 Midori_U381 ( .A(wk_share3[6]), .B(Midori_rounds_SR_Result3[46]), 
        .Z(output3[6]) );
  XOR2_X1 Midori_U380 ( .A(wk_share3[63]), .B(Midori_rounds_SR_Result3[63]), 
        .Z(output3[63]) );
  XOR2_X1 Midori_U379 ( .A(wk_share3[62]), .B(Midori_rounds_SR_Result3[62]), 
        .Z(output3[62]) );
  XOR2_X1 Midori_U378 ( .A(wk_share3[61]), .B(Midori_rounds_SR_Result3[61]), 
        .Z(output3[61]) );
  XOR2_X1 Midori_U377 ( .A(wk_share3[60]), .B(Midori_rounds_SR_Result3[60]), 
        .Z(output3[60]) );
  XOR2_X1 Midori_U376 ( .A(wk_share3[5]), .B(Midori_rounds_SR_Result3[45]), 
        .Z(output3[5]) );
  XOR2_X1 Midori_U375 ( .A(wk_share3[59]), .B(Midori_rounds_SR_Result3[35]), 
        .Z(output3[59]) );
  XOR2_X1 Midori_U374 ( .A(wk_share3[58]), .B(Midori_rounds_SR_Result3[34]), 
        .Z(output3[58]) );
  XOR2_X1 Midori_U373 ( .A(wk_share3[57]), .B(Midori_rounds_SR_Result3[33]), 
        .Z(output3[57]) );
  XOR2_X1 Midori_U372 ( .A(wk_share3[56]), .B(Midori_rounds_SR_Result3[32]), 
        .Z(output3[56]) );
  XOR2_X1 Midori_U371 ( .A(wk_share3[55]), .B(Midori_rounds_SR_Result3[7]), 
        .Z(output3[55]) );
  XOR2_X1 Midori_U370 ( .A(wk_share3[54]), .B(Midori_rounds_SR_Result3[6]), 
        .Z(output3[54]) );
  XOR2_X1 Midori_U369 ( .A(wk_share3[53]), .B(Midori_rounds_SR_Result3[5]), 
        .Z(output3[53]) );
  XOR2_X1 Midori_U368 ( .A(wk_share3[52]), .B(Midori_rounds_SR_Result3[4]), 
        .Z(output3[52]) );
  XOR2_X1 Midori_U367 ( .A(wk_share3[51]), .B(Midori_rounds_SR_Result3[27]), 
        .Z(output3[51]) );
  XOR2_X1 Midori_U366 ( .A(wk_share3[50]), .B(Midori_rounds_SR_Result3[26]), 
        .Z(output3[50]) );
  XOR2_X1 Midori_U365 ( .A(wk_share3[4]), .B(Midori_rounds_SR_Result3[44]), 
        .Z(output3[4]) );
  XOR2_X1 Midori_U364 ( .A(wk_share3[49]), .B(Midori_rounds_SR_Result3[25]), 
        .Z(output3[49]) );
  XOR2_X1 Midori_U363 ( .A(wk_share3[48]), .B(Midori_rounds_SR_Result3[24]), 
        .Z(output3[48]) );
  XOR2_X1 Midori_U362 ( .A(wk_share3[47]), .B(Midori_rounds_SR_Result3[43]), 
        .Z(output3[47]) );
  XOR2_X1 Midori_U361 ( .A(wk_share3[46]), .B(Midori_rounds_SR_Result3[42]), 
        .Z(output3[46]) );
  XOR2_X1 Midori_U360 ( .A(wk_share3[45]), .B(Midori_rounds_SR_Result3[41]), 
        .Z(output3[45]) );
  XOR2_X1 Midori_U359 ( .A(wk_share3[44]), .B(Midori_rounds_SR_Result3[40]), 
        .Z(output3[44]) );
  XOR2_X1 Midori_U358 ( .A(wk_share3[43]), .B(Midori_rounds_SR_Result3[55]), 
        .Z(output3[43]) );
  XOR2_X1 Midori_U357 ( .A(wk_share3[42]), .B(Midori_rounds_SR_Result3[54]), 
        .Z(output3[42]) );
  XOR2_X1 Midori_U356 ( .A(wk_share3[41]), .B(Midori_rounds_SR_Result3[53]), 
        .Z(output3[41]) );
  XOR2_X1 Midori_U355 ( .A(wk_share3[40]), .B(Midori_rounds_SR_Result3[52]), 
        .Z(output3[40]) );
  XOR2_X1 Midori_U354 ( .A(wk_share3[3]), .B(Midori_rounds_SR_Result3[51]), 
        .Z(output3[3]) );
  XOR2_X1 Midori_U353 ( .A(wk_share3[39]), .B(Midori_rounds_SR_Result3[19]), 
        .Z(output3[39]) );
  XOR2_X1 Midori_U352 ( .A(wk_share3[38]), .B(Midori_rounds_SR_Result3[18]), 
        .Z(output3[38]) );
  XOR2_X1 Midori_U351 ( .A(wk_share3[37]), .B(Midori_rounds_SR_Result3[17]), 
        .Z(output3[37]) );
  XOR2_X1 Midori_U350 ( .A(wk_share3[36]), .B(Midori_rounds_SR_Result3[16]), 
        .Z(output3[36]) );
  XOR2_X1 Midori_U349 ( .A(wk_share3[35]), .B(Midori_rounds_SR_Result3[15]), 
        .Z(output3[35]) );
  XOR2_X1 Midori_U348 ( .A(wk_share3[34]), .B(Midori_rounds_SR_Result3[14]), 
        .Z(output3[34]) );
  XOR2_X1 Midori_U347 ( .A(wk_share3[33]), .B(Midori_rounds_SR_Result3[13]), 
        .Z(output3[33]) );
  XOR2_X1 Midori_U346 ( .A(wk_share3[32]), .B(Midori_rounds_SR_Result3[12]), 
        .Z(output3[32]) );
  XOR2_X1 Midori_U345 ( .A(wk_share3[31]), .B(Midori_rounds_SR_Result3[3]), 
        .Z(output3[31]) );
  XOR2_X1 Midori_U344 ( .A(wk_share3[30]), .B(Midori_rounds_SR_Result3[2]), 
        .Z(output3[30]) );
  XOR2_X1 Midori_U343 ( .A(wk_share3[2]), .B(Midori_rounds_SR_Result3[50]), 
        .Z(output3[2]) );
  XOR2_X1 Midori_U342 ( .A(wk_share3[29]), .B(Midori_rounds_SR_Result3[1]), 
        .Z(output3[29]) );
  XOR2_X1 Midori_U341 ( .A(wk_share3[28]), .B(Midori_rounds_SR_Result3[0]), 
        .Z(output3[28]) );
  XOR2_X1 Midori_U340 ( .A(wk_share3[27]), .B(Midori_rounds_SR_Result3[31]), 
        .Z(output3[27]) );
  XOR2_X1 Midori_U339 ( .A(wk_share3[26]), .B(Midori_rounds_SR_Result3[30]), 
        .Z(output3[26]) );
  XOR2_X1 Midori_U338 ( .A(wk_share3[25]), .B(Midori_rounds_SR_Result3[29]), 
        .Z(output3[25]) );
  XOR2_X1 Midori_U337 ( .A(wk_share3[24]), .B(Midori_rounds_SR_Result3[28]), 
        .Z(output3[24]) );
  XOR2_X1 Midori_U336 ( .A(wk_share3[23]), .B(Midori_rounds_SR_Result3[59]), 
        .Z(output3[23]) );
  XOR2_X1 Midori_U335 ( .A(wk_share3[22]), .B(Midori_rounds_SR_Result3[58]), 
        .Z(output3[22]) );
  XOR2_X1 Midori_U334 ( .A(wk_share3[21]), .B(Midori_rounds_SR_Result3[57]), 
        .Z(output3[21]) );
  XOR2_X1 Midori_U333 ( .A(wk_share3[20]), .B(Midori_rounds_SR_Result3[56]), 
        .Z(output3[20]) );
  XOR2_X1 Midori_U332 ( .A(wk_share3[1]), .B(Midori_rounds_SR_Result3[49]), 
        .Z(output3[1]) );
  XOR2_X1 Midori_U331 ( .A(wk_share3[19]), .B(Midori_rounds_SR_Result3[39]), 
        .Z(output3[19]) );
  XOR2_X1 Midori_U330 ( .A(wk_share3[18]), .B(Midori_rounds_SR_Result3[38]), 
        .Z(output3[18]) );
  XOR2_X1 Midori_U329 ( .A(wk_share3[17]), .B(Midori_rounds_SR_Result3[37]), 
        .Z(output3[17]) );
  XOR2_X1 Midori_U328 ( .A(wk_share3[16]), .B(Midori_rounds_SR_Result3[36]), 
        .Z(output3[16]) );
  XOR2_X1 Midori_U327 ( .A(wk_share3[15]), .B(Midori_rounds_SR_Result3[23]), 
        .Z(output3[15]) );
  XOR2_X1 Midori_U326 ( .A(wk_share3[14]), .B(Midori_rounds_SR_Result3[22]), 
        .Z(output3[14]) );
  XOR2_X1 Midori_U325 ( .A(wk_share3[13]), .B(Midori_rounds_SR_Result3[21]), 
        .Z(output3[13]) );
  XOR2_X1 Midori_U324 ( .A(wk_share3[12]), .B(Midori_rounds_SR_Result3[20]), 
        .Z(output3[12]) );
  XOR2_X1 Midori_U323 ( .A(wk_share3[11]), .B(Midori_rounds_SR_Result3[11]), 
        .Z(output3[11]) );
  XOR2_X1 Midori_U322 ( .A(wk_share3[10]), .B(Midori_rounds_SR_Result3[10]), 
        .Z(output3[10]) );
  XOR2_X1 Midori_U321 ( .A(wk_share3[0]), .B(Midori_rounds_SR_Result3[48]), 
        .Z(output3[0]) );
  XOR2_X1 Midori_U320 ( .A(wk_share2[9]), .B(Midori_rounds_SR_Result2[9]), .Z(
        output2[9]) );
  XOR2_X1 Midori_U319 ( .A(wk_share2[8]), .B(Midori_rounds_SR_Result2[8]), .Z(
        output2[8]) );
  XOR2_X1 Midori_U318 ( .A(wk_share2[7]), .B(Midori_rounds_SR_Result2[47]), 
        .Z(output2[7]) );
  XOR2_X1 Midori_U317 ( .A(wk_share2[6]), .B(Midori_rounds_SR_Result2[46]), 
        .Z(output2[6]) );
  XOR2_X1 Midori_U316 ( .A(wk_share2[63]), .B(Midori_rounds_SR_Result2[63]), 
        .Z(output2[63]) );
  XOR2_X1 Midori_U315 ( .A(wk_share2[62]), .B(Midori_rounds_SR_Result2[62]), 
        .Z(output2[62]) );
  XOR2_X1 Midori_U314 ( .A(wk_share2[61]), .B(Midori_rounds_SR_Result2[61]), 
        .Z(output2[61]) );
  XOR2_X1 Midori_U313 ( .A(wk_share2[60]), .B(Midori_rounds_SR_Result2[60]), 
        .Z(output2[60]) );
  XOR2_X1 Midori_U312 ( .A(wk_share2[5]), .B(Midori_rounds_SR_Result2[45]), 
        .Z(output2[5]) );
  XOR2_X1 Midori_U311 ( .A(wk_share2[59]), .B(Midori_rounds_SR_Result2[35]), 
        .Z(output2[59]) );
  XOR2_X1 Midori_U310 ( .A(wk_share2[58]), .B(Midori_rounds_SR_Result2[34]), 
        .Z(output2[58]) );
  XOR2_X1 Midori_U309 ( .A(wk_share2[57]), .B(Midori_rounds_SR_Result2[33]), 
        .Z(output2[57]) );
  XOR2_X1 Midori_U308 ( .A(wk_share2[56]), .B(Midori_rounds_SR_Result2[32]), 
        .Z(output2[56]) );
  XOR2_X1 Midori_U307 ( .A(wk_share2[55]), .B(Midori_rounds_SR_Result2[7]), 
        .Z(output2[55]) );
  XOR2_X1 Midori_U306 ( .A(wk_share2[54]), .B(Midori_rounds_SR_Result2[6]), 
        .Z(output2[54]) );
  XOR2_X1 Midori_U305 ( .A(wk_share2[53]), .B(Midori_rounds_SR_Result2[5]), 
        .Z(output2[53]) );
  XOR2_X1 Midori_U304 ( .A(wk_share2[52]), .B(Midori_rounds_SR_Result2[4]), 
        .Z(output2[52]) );
  XOR2_X1 Midori_U303 ( .A(wk_share2[51]), .B(Midori_rounds_SR_Result2[27]), 
        .Z(output2[51]) );
  XOR2_X1 Midori_U302 ( .A(wk_share2[50]), .B(Midori_rounds_SR_Result2[26]), 
        .Z(output2[50]) );
  XOR2_X1 Midori_U301 ( .A(wk_share2[4]), .B(Midori_rounds_SR_Result2[44]), 
        .Z(output2[4]) );
  XOR2_X1 Midori_U300 ( .A(wk_share2[49]), .B(Midori_rounds_SR_Result2[25]), 
        .Z(output2[49]) );
  XOR2_X1 Midori_U299 ( .A(wk_share2[48]), .B(Midori_rounds_SR_Result2[24]), 
        .Z(output2[48]) );
  XOR2_X1 Midori_U298 ( .A(wk_share2[47]), .B(Midori_rounds_SR_Result2[43]), 
        .Z(output2[47]) );
  XOR2_X1 Midori_U297 ( .A(wk_share2[46]), .B(Midori_rounds_SR_Result2[42]), 
        .Z(output2[46]) );
  XOR2_X1 Midori_U296 ( .A(wk_share2[45]), .B(Midori_rounds_SR_Result2[41]), 
        .Z(output2[45]) );
  XOR2_X1 Midori_U295 ( .A(wk_share2[44]), .B(Midori_rounds_SR_Result2[40]), 
        .Z(output2[44]) );
  XOR2_X1 Midori_U294 ( .A(wk_share2[43]), .B(Midori_rounds_SR_Result2[55]), 
        .Z(output2[43]) );
  XOR2_X1 Midori_U293 ( .A(wk_share2[42]), .B(Midori_rounds_SR_Result2[54]), 
        .Z(output2[42]) );
  XOR2_X1 Midori_U292 ( .A(wk_share2[41]), .B(Midori_rounds_SR_Result2[53]), 
        .Z(output2[41]) );
  XOR2_X1 Midori_U291 ( .A(wk_share2[40]), .B(Midori_rounds_SR_Result2[52]), 
        .Z(output2[40]) );
  XOR2_X1 Midori_U290 ( .A(wk_share2[3]), .B(Midori_rounds_SR_Result2[51]), 
        .Z(output2[3]) );
  XOR2_X1 Midori_U289 ( .A(wk_share2[39]), .B(Midori_rounds_SR_Result2[19]), 
        .Z(output2[39]) );
  XOR2_X1 Midori_U288 ( .A(wk_share2[38]), .B(Midori_rounds_SR_Result2[18]), 
        .Z(output2[38]) );
  XOR2_X1 Midori_U287 ( .A(wk_share2[37]), .B(Midori_rounds_SR_Result2[17]), 
        .Z(output2[37]) );
  XOR2_X1 Midori_U286 ( .A(wk_share2[36]), .B(Midori_rounds_SR_Result2[16]), 
        .Z(output2[36]) );
  XOR2_X1 Midori_U285 ( .A(wk_share2[35]), .B(Midori_rounds_SR_Result2[15]), 
        .Z(output2[35]) );
  XOR2_X1 Midori_U284 ( .A(wk_share2[34]), .B(Midori_rounds_SR_Result2[14]), 
        .Z(output2[34]) );
  XOR2_X1 Midori_U283 ( .A(wk_share2[33]), .B(Midori_rounds_SR_Result2[13]), 
        .Z(output2[33]) );
  XOR2_X1 Midori_U282 ( .A(wk_share2[32]), .B(Midori_rounds_SR_Result2[12]), 
        .Z(output2[32]) );
  XOR2_X1 Midori_U281 ( .A(wk_share2[31]), .B(Midori_rounds_SR_Result2[3]), 
        .Z(output2[31]) );
  XOR2_X1 Midori_U280 ( .A(wk_share2[30]), .B(Midori_rounds_SR_Result2[2]), 
        .Z(output2[30]) );
  XOR2_X1 Midori_U279 ( .A(wk_share2[2]), .B(Midori_rounds_SR_Result2[50]), 
        .Z(output2[2]) );
  XOR2_X1 Midori_U278 ( .A(wk_share2[29]), .B(Midori_rounds_SR_Result2[1]), 
        .Z(output2[29]) );
  XOR2_X1 Midori_U277 ( .A(wk_share2[28]), .B(Midori_rounds_SR_Result2[0]), 
        .Z(output2[28]) );
  XOR2_X1 Midori_U276 ( .A(wk_share2[27]), .B(Midori_rounds_SR_Result2[31]), 
        .Z(output2[27]) );
  XOR2_X1 Midori_U275 ( .A(wk_share2[26]), .B(Midori_rounds_SR_Result2[30]), 
        .Z(output2[26]) );
  XOR2_X1 Midori_U274 ( .A(wk_share2[25]), .B(Midori_rounds_SR_Result2[29]), 
        .Z(output2[25]) );
  XOR2_X1 Midori_U273 ( .A(wk_share2[24]), .B(Midori_rounds_SR_Result2[28]), 
        .Z(output2[24]) );
  XOR2_X1 Midori_U272 ( .A(wk_share2[23]), .B(Midori_rounds_SR_Result2[59]), 
        .Z(output2[23]) );
  XOR2_X1 Midori_U271 ( .A(wk_share2[22]), .B(Midori_rounds_SR_Result2[58]), 
        .Z(output2[22]) );
  XOR2_X1 Midori_U270 ( .A(wk_share2[21]), .B(Midori_rounds_SR_Result2[57]), 
        .Z(output2[21]) );
  XOR2_X1 Midori_U269 ( .A(wk_share2[20]), .B(Midori_rounds_SR_Result2[56]), 
        .Z(output2[20]) );
  XOR2_X1 Midori_U268 ( .A(wk_share2[1]), .B(Midori_rounds_SR_Result2[49]), 
        .Z(output2[1]) );
  XOR2_X1 Midori_U267 ( .A(wk_share2[19]), .B(Midori_rounds_SR_Result2[39]), 
        .Z(output2[19]) );
  XOR2_X1 Midori_U266 ( .A(wk_share2[18]), .B(Midori_rounds_SR_Result2[38]), 
        .Z(output2[18]) );
  XOR2_X1 Midori_U265 ( .A(wk_share2[17]), .B(Midori_rounds_SR_Result2[37]), 
        .Z(output2[17]) );
  XOR2_X1 Midori_U264 ( .A(wk_share2[16]), .B(Midori_rounds_SR_Result2[36]), 
        .Z(output2[16]) );
  XOR2_X1 Midori_U263 ( .A(wk_share2[15]), .B(Midori_rounds_SR_Result2[23]), 
        .Z(output2[15]) );
  XOR2_X1 Midori_U262 ( .A(wk_share2[14]), .B(Midori_rounds_SR_Result2[22]), 
        .Z(output2[14]) );
  XOR2_X1 Midori_U261 ( .A(wk_share2[13]), .B(Midori_rounds_SR_Result2[21]), 
        .Z(output2[13]) );
  XOR2_X1 Midori_U260 ( .A(wk_share2[12]), .B(Midori_rounds_SR_Result2[20]), 
        .Z(output2[12]) );
  XOR2_X1 Midori_U259 ( .A(wk_share2[11]), .B(Midori_rounds_SR_Result2[11]), 
        .Z(output2[11]) );
  XOR2_X1 Midori_U258 ( .A(wk_share2[10]), .B(Midori_rounds_SR_Result2[10]), 
        .Z(output2[10]) );
  XOR2_X1 Midori_U257 ( .A(wk_share2[0]), .B(Midori_rounds_SR_Result2[48]), 
        .Z(output2[0]) );
  XOR2_X1 Midori_U256 ( .A(wk_share1[9]), .B(Midori_rounds_SR_Result1[9]), .Z(
        output1[9]) );
  XOR2_X1 Midori_U255 ( .A(wk_share1[8]), .B(Midori_rounds_SR_Result1[8]), .Z(
        output1[8]) );
  XOR2_X1 Midori_U254 ( .A(wk_share1[7]), .B(Midori_rounds_SR_Result1[47]), 
        .Z(output1[7]) );
  XOR2_X1 Midori_U253 ( .A(wk_share1[6]), .B(Midori_rounds_SR_Result1[46]), 
        .Z(output1[6]) );
  XOR2_X1 Midori_U252 ( .A(wk_share1[63]), .B(Midori_rounds_SR_Result1[63]), 
        .Z(output1[63]) );
  XOR2_X1 Midori_U251 ( .A(wk_share1[62]), .B(Midori_rounds_SR_Result1[62]), 
        .Z(output1[62]) );
  XOR2_X1 Midori_U250 ( .A(wk_share1[61]), .B(Midori_rounds_SR_Result1[61]), 
        .Z(output1[61]) );
  XOR2_X1 Midori_U249 ( .A(wk_share1[60]), .B(Midori_rounds_SR_Result1[60]), 
        .Z(output1[60]) );
  XOR2_X1 Midori_U248 ( .A(wk_share1[5]), .B(Midori_rounds_SR_Result1[45]), 
        .Z(output1[5]) );
  XOR2_X1 Midori_U247 ( .A(wk_share1[59]), .B(Midori_rounds_SR_Result1[35]), 
        .Z(output1[59]) );
  XOR2_X1 Midori_U246 ( .A(wk_share1[58]), .B(Midori_rounds_SR_Result1[34]), 
        .Z(output1[58]) );
  XOR2_X1 Midori_U245 ( .A(wk_share1[57]), .B(Midori_rounds_SR_Result1[33]), 
        .Z(output1[57]) );
  XOR2_X1 Midori_U244 ( .A(wk_share1[56]), .B(Midori_rounds_SR_Result1[32]), 
        .Z(output1[56]) );
  XOR2_X1 Midori_U243 ( .A(wk_share1[55]), .B(Midori_rounds_SR_Result1[7]), 
        .Z(output1[55]) );
  XOR2_X1 Midori_U242 ( .A(wk_share1[54]), .B(Midori_rounds_SR_Result1[6]), 
        .Z(output1[54]) );
  XOR2_X1 Midori_U241 ( .A(wk_share1[53]), .B(Midori_rounds_SR_Result1[5]), 
        .Z(output1[53]) );
  XOR2_X1 Midori_U240 ( .A(wk_share1[52]), .B(Midori_rounds_SR_Result1[4]), 
        .Z(output1[52]) );
  XOR2_X1 Midori_U239 ( .A(wk_share1[51]), .B(Midori_rounds_SR_Result1[27]), 
        .Z(output1[51]) );
  XOR2_X1 Midori_U238 ( .A(wk_share1[50]), .B(Midori_rounds_SR_Result1[26]), 
        .Z(output1[50]) );
  XOR2_X1 Midori_U237 ( .A(wk_share1[4]), .B(Midori_rounds_SR_Result1[44]), 
        .Z(output1[4]) );
  XOR2_X1 Midori_U236 ( .A(wk_share1[49]), .B(Midori_rounds_SR_Result1[25]), 
        .Z(output1[49]) );
  XOR2_X1 Midori_U235 ( .A(wk_share1[48]), .B(Midori_rounds_SR_Result1[24]), 
        .Z(output1[48]) );
  XOR2_X1 Midori_U234 ( .A(wk_share1[47]), .B(Midori_rounds_SR_Result1[43]), 
        .Z(output1[47]) );
  XOR2_X1 Midori_U233 ( .A(wk_share1[46]), .B(Midori_rounds_SR_Result1[42]), 
        .Z(output1[46]) );
  XOR2_X1 Midori_U232 ( .A(wk_share1[45]), .B(Midori_rounds_SR_Result1[41]), 
        .Z(output1[45]) );
  XOR2_X1 Midori_U231 ( .A(wk_share1[44]), .B(Midori_rounds_SR_Result1[40]), 
        .Z(output1[44]) );
  XOR2_X1 Midori_U230 ( .A(wk_share1[43]), .B(Midori_rounds_SR_Result1[55]), 
        .Z(output1[43]) );
  XOR2_X1 Midori_U229 ( .A(wk_share1[42]), .B(Midori_rounds_SR_Result1[54]), 
        .Z(output1[42]) );
  XOR2_X1 Midori_U228 ( .A(wk_share1[41]), .B(Midori_rounds_SR_Result1[53]), 
        .Z(output1[41]) );
  XOR2_X1 Midori_U227 ( .A(wk_share1[40]), .B(Midori_rounds_SR_Result1[52]), 
        .Z(output1[40]) );
  XOR2_X1 Midori_U226 ( .A(wk_share1[3]), .B(Midori_rounds_SR_Result1[51]), 
        .Z(output1[3]) );
  XOR2_X1 Midori_U225 ( .A(wk_share1[39]), .B(Midori_rounds_SR_Result1[19]), 
        .Z(output1[39]) );
  XOR2_X1 Midori_U224 ( .A(wk_share1[38]), .B(Midori_rounds_SR_Result1[18]), 
        .Z(output1[38]) );
  XOR2_X1 Midori_U223 ( .A(wk_share1[37]), .B(Midori_rounds_SR_Result1[17]), 
        .Z(output1[37]) );
  XOR2_X1 Midori_U222 ( .A(wk_share1[36]), .B(Midori_rounds_SR_Result1[16]), 
        .Z(output1[36]) );
  XOR2_X1 Midori_U221 ( .A(wk_share1[35]), .B(Midori_rounds_SR_Result1[15]), 
        .Z(output1[35]) );
  XOR2_X1 Midori_U220 ( .A(wk_share1[34]), .B(Midori_rounds_SR_Result1[14]), 
        .Z(output1[34]) );
  XOR2_X1 Midori_U219 ( .A(wk_share1[33]), .B(Midori_rounds_SR_Result1[13]), 
        .Z(output1[33]) );
  XOR2_X1 Midori_U218 ( .A(wk_share1[32]), .B(Midori_rounds_SR_Result1[12]), 
        .Z(output1[32]) );
  XOR2_X1 Midori_U217 ( .A(wk_share1[31]), .B(Midori_rounds_SR_Result1[3]), 
        .Z(output1[31]) );
  XOR2_X1 Midori_U216 ( .A(wk_share1[30]), .B(Midori_rounds_SR_Result1[2]), 
        .Z(output1[30]) );
  XOR2_X1 Midori_U215 ( .A(wk_share1[2]), .B(Midori_rounds_SR_Result1[50]), 
        .Z(output1[2]) );
  XOR2_X1 Midori_U214 ( .A(wk_share1[29]), .B(Midori_rounds_SR_Result1[1]), 
        .Z(output1[29]) );
  XOR2_X1 Midori_U213 ( .A(wk_share1[28]), .B(Midori_rounds_SR_Result1[0]), 
        .Z(output1[28]) );
  XOR2_X1 Midori_U212 ( .A(wk_share1[27]), .B(Midori_rounds_SR_Result1[31]), 
        .Z(output1[27]) );
  XOR2_X1 Midori_U211 ( .A(wk_share1[26]), .B(Midori_rounds_SR_Result1[30]), 
        .Z(output1[26]) );
  XOR2_X1 Midori_U210 ( .A(wk_share1[25]), .B(Midori_rounds_SR_Result1[29]), 
        .Z(output1[25]) );
  XOR2_X1 Midori_U209 ( .A(wk_share1[24]), .B(Midori_rounds_SR_Result1[28]), 
        .Z(output1[24]) );
  XOR2_X1 Midori_U208 ( .A(wk_share1[23]), .B(Midori_rounds_SR_Result1[59]), 
        .Z(output1[23]) );
  XOR2_X1 Midori_U207 ( .A(wk_share1[22]), .B(Midori_rounds_SR_Result1[58]), 
        .Z(output1[22]) );
  XOR2_X1 Midori_U206 ( .A(wk_share1[21]), .B(Midori_rounds_SR_Result1[57]), 
        .Z(output1[21]) );
  XOR2_X1 Midori_U205 ( .A(wk_share1[20]), .B(Midori_rounds_SR_Result1[56]), 
        .Z(output1[20]) );
  XOR2_X1 Midori_U204 ( .A(wk_share1[1]), .B(Midori_rounds_SR_Result1[49]), 
        .Z(output1[1]) );
  XOR2_X1 Midori_U203 ( .A(wk_share1[19]), .B(Midori_rounds_SR_Result1[39]), 
        .Z(output1[19]) );
  XOR2_X1 Midori_U202 ( .A(wk_share1[18]), .B(Midori_rounds_SR_Result1[38]), 
        .Z(output1[18]) );
  XOR2_X1 Midori_U201 ( .A(wk_share1[17]), .B(Midori_rounds_SR_Result1[37]), 
        .Z(output1[17]) );
  XOR2_X1 Midori_U200 ( .A(wk_share1[16]), .B(Midori_rounds_SR_Result1[36]), 
        .Z(output1[16]) );
  XOR2_X1 Midori_U199 ( .A(wk_share1[15]), .B(Midori_rounds_SR_Result1[23]), 
        .Z(output1[15]) );
  XOR2_X1 Midori_U198 ( .A(wk_share1[14]), .B(Midori_rounds_SR_Result1[22]), 
        .Z(output1[14]) );
  XOR2_X1 Midori_U197 ( .A(wk_share1[13]), .B(Midori_rounds_SR_Result1[21]), 
        .Z(output1[13]) );
  XOR2_X1 Midori_U196 ( .A(wk_share1[12]), .B(Midori_rounds_SR_Result1[20]), 
        .Z(output1[12]) );
  XOR2_X1 Midori_U195 ( .A(wk_share1[11]), .B(Midori_rounds_SR_Result1[11]), 
        .Z(output1[11]) );
  XOR2_X1 Midori_U194 ( .A(wk_share1[10]), .B(Midori_rounds_SR_Result1[10]), 
        .Z(output1[10]) );
  XOR2_X1 Midori_U193 ( .A(wk_share1[0]), .B(Midori_rounds_SR_Result1[48]), 
        .Z(output1[0]) );
  XOR2_X1 Midori_U192 ( .A(wk_share3[9]), .B(input3[9]), .Z(
        Midori_add_Result_Start3[9]) );
  XOR2_X1 Midori_U191 ( .A(wk_share3[8]), .B(input3[8]), .Z(
        Midori_add_Result_Start3[8]) );
  XOR2_X1 Midori_U190 ( .A(wk_share3[7]), .B(input3[7]), .Z(
        Midori_add_Result_Start3[7]) );
  XOR2_X1 Midori_U189 ( .A(wk_share3[6]), .B(input3[6]), .Z(
        Midori_add_Result_Start3[6]) );
  XOR2_X1 Midori_U188 ( .A(wk_share3[63]), .B(input3[63]), .Z(
        Midori_add_Result_Start3[63]) );
  XOR2_X1 Midori_U187 ( .A(wk_share3[62]), .B(input3[62]), .Z(
        Midori_add_Result_Start3[62]) );
  XOR2_X1 Midori_U186 ( .A(wk_share3[61]), .B(input3[61]), .Z(
        Midori_add_Result_Start3[61]) );
  XOR2_X1 Midori_U185 ( .A(wk_share3[60]), .B(input3[60]), .Z(
        Midori_add_Result_Start3[60]) );
  XOR2_X1 Midori_U184 ( .A(wk_share3[5]), .B(input3[5]), .Z(
        Midori_add_Result_Start3[5]) );
  XOR2_X1 Midori_U183 ( .A(wk_share3[59]), .B(input3[59]), .Z(
        Midori_add_Result_Start3[59]) );
  XOR2_X1 Midori_U182 ( .A(wk_share3[58]), .B(input3[58]), .Z(
        Midori_add_Result_Start3[58]) );
  XOR2_X1 Midori_U181 ( .A(wk_share3[57]), .B(input3[57]), .Z(
        Midori_add_Result_Start3[57]) );
  XOR2_X1 Midori_U180 ( .A(wk_share3[56]), .B(input3[56]), .Z(
        Midori_add_Result_Start3[56]) );
  XOR2_X1 Midori_U179 ( .A(wk_share3[55]), .B(input3[55]), .Z(
        Midori_add_Result_Start3[55]) );
  XOR2_X1 Midori_U178 ( .A(wk_share3[54]), .B(input3[54]), .Z(
        Midori_add_Result_Start3[54]) );
  XOR2_X1 Midori_U177 ( .A(wk_share3[53]), .B(input3[53]), .Z(
        Midori_add_Result_Start3[53]) );
  XOR2_X1 Midori_U176 ( .A(wk_share3[52]), .B(input3[52]), .Z(
        Midori_add_Result_Start3[52]) );
  XOR2_X1 Midori_U175 ( .A(wk_share3[51]), .B(input3[51]), .Z(
        Midori_add_Result_Start3[51]) );
  XOR2_X1 Midori_U174 ( .A(wk_share3[50]), .B(input3[50]), .Z(
        Midori_add_Result_Start3[50]) );
  XOR2_X1 Midori_U173 ( .A(wk_share3[4]), .B(input3[4]), .Z(
        Midori_add_Result_Start3[4]) );
  XOR2_X1 Midori_U172 ( .A(wk_share3[49]), .B(input3[49]), .Z(
        Midori_add_Result_Start3[49]) );
  XOR2_X1 Midori_U171 ( .A(wk_share3[48]), .B(input3[48]), .Z(
        Midori_add_Result_Start3[48]) );
  XOR2_X1 Midori_U170 ( .A(wk_share3[47]), .B(input3[47]), .Z(
        Midori_add_Result_Start3[47]) );
  XOR2_X1 Midori_U169 ( .A(wk_share3[46]), .B(input3[46]), .Z(
        Midori_add_Result_Start3[46]) );
  XOR2_X1 Midori_U168 ( .A(wk_share3[45]), .B(input3[45]), .Z(
        Midori_add_Result_Start3[45]) );
  XOR2_X1 Midori_U167 ( .A(wk_share3[44]), .B(input3[44]), .Z(
        Midori_add_Result_Start3[44]) );
  XOR2_X1 Midori_U166 ( .A(wk_share3[43]), .B(input3[43]), .Z(
        Midori_add_Result_Start3[43]) );
  XOR2_X1 Midori_U165 ( .A(wk_share3[42]), .B(input3[42]), .Z(
        Midori_add_Result_Start3[42]) );
  XOR2_X1 Midori_U164 ( .A(wk_share3[41]), .B(input3[41]), .Z(
        Midori_add_Result_Start3[41]) );
  XOR2_X1 Midori_U163 ( .A(wk_share3[40]), .B(input3[40]), .Z(
        Midori_add_Result_Start3[40]) );
  XOR2_X1 Midori_U162 ( .A(wk_share3[3]), .B(input3[3]), .Z(
        Midori_add_Result_Start3[3]) );
  XOR2_X1 Midori_U161 ( .A(wk_share3[39]), .B(input3[39]), .Z(
        Midori_add_Result_Start3[39]) );
  XOR2_X1 Midori_U160 ( .A(wk_share3[38]), .B(input3[38]), .Z(
        Midori_add_Result_Start3[38]) );
  XOR2_X1 Midori_U159 ( .A(wk_share3[37]), .B(input3[37]), .Z(
        Midori_add_Result_Start3[37]) );
  XOR2_X1 Midori_U158 ( .A(wk_share3[36]), .B(input3[36]), .Z(
        Midori_add_Result_Start3[36]) );
  XOR2_X1 Midori_U157 ( .A(wk_share3[35]), .B(input3[35]), .Z(
        Midori_add_Result_Start3[35]) );
  XOR2_X1 Midori_U156 ( .A(wk_share3[34]), .B(input3[34]), .Z(
        Midori_add_Result_Start3[34]) );
  XOR2_X1 Midori_U155 ( .A(wk_share3[33]), .B(input3[33]), .Z(
        Midori_add_Result_Start3[33]) );
  XOR2_X1 Midori_U154 ( .A(wk_share3[32]), .B(input3[32]), .Z(
        Midori_add_Result_Start3[32]) );
  XOR2_X1 Midori_U153 ( .A(wk_share3[31]), .B(input3[31]), .Z(
        Midori_add_Result_Start3[31]) );
  XOR2_X1 Midori_U152 ( .A(wk_share3[30]), .B(input3[30]), .Z(
        Midori_add_Result_Start3[30]) );
  XOR2_X1 Midori_U151 ( .A(wk_share3[2]), .B(input3[2]), .Z(
        Midori_add_Result_Start3[2]) );
  XOR2_X1 Midori_U150 ( .A(wk_share3[29]), .B(input3[29]), .Z(
        Midori_add_Result_Start3[29]) );
  XOR2_X1 Midori_U149 ( .A(wk_share3[28]), .B(input3[28]), .Z(
        Midori_add_Result_Start3[28]) );
  XOR2_X1 Midori_U148 ( .A(wk_share3[27]), .B(input3[27]), .Z(
        Midori_add_Result_Start3[27]) );
  XOR2_X1 Midori_U147 ( .A(wk_share3[26]), .B(input3[26]), .Z(
        Midori_add_Result_Start3[26]) );
  XOR2_X1 Midori_U146 ( .A(wk_share3[25]), .B(input3[25]), .Z(
        Midori_add_Result_Start3[25]) );
  XOR2_X1 Midori_U145 ( .A(wk_share3[24]), .B(input3[24]), .Z(
        Midori_add_Result_Start3[24]) );
  XOR2_X1 Midori_U144 ( .A(wk_share3[23]), .B(input3[23]), .Z(
        Midori_add_Result_Start3[23]) );
  XOR2_X1 Midori_U143 ( .A(wk_share3[22]), .B(input3[22]), .Z(
        Midori_add_Result_Start3[22]) );
  XOR2_X1 Midori_U142 ( .A(wk_share3[21]), .B(input3[21]), .Z(
        Midori_add_Result_Start3[21]) );
  XOR2_X1 Midori_U141 ( .A(wk_share3[20]), .B(input3[20]), .Z(
        Midori_add_Result_Start3[20]) );
  XOR2_X1 Midori_U140 ( .A(wk_share3[1]), .B(input3[1]), .Z(
        Midori_add_Result_Start3[1]) );
  XOR2_X1 Midori_U139 ( .A(wk_share3[19]), .B(input3[19]), .Z(
        Midori_add_Result_Start3[19]) );
  XOR2_X1 Midori_U138 ( .A(wk_share3[18]), .B(input3[18]), .Z(
        Midori_add_Result_Start3[18]) );
  XOR2_X1 Midori_U137 ( .A(wk_share3[17]), .B(input3[17]), .Z(
        Midori_add_Result_Start3[17]) );
  XOR2_X1 Midori_U136 ( .A(wk_share3[16]), .B(input3[16]), .Z(
        Midori_add_Result_Start3[16]) );
  XOR2_X1 Midori_U135 ( .A(wk_share3[15]), .B(input3[15]), .Z(
        Midori_add_Result_Start3[15]) );
  XOR2_X1 Midori_U134 ( .A(wk_share3[14]), .B(input3[14]), .Z(
        Midori_add_Result_Start3[14]) );
  XOR2_X1 Midori_U133 ( .A(wk_share3[13]), .B(input3[13]), .Z(
        Midori_add_Result_Start3[13]) );
  XOR2_X1 Midori_U132 ( .A(wk_share3[12]), .B(input3[12]), .Z(
        Midori_add_Result_Start3[12]) );
  XOR2_X1 Midori_U131 ( .A(wk_share3[11]), .B(input3[11]), .Z(
        Midori_add_Result_Start3[11]) );
  XOR2_X1 Midori_U130 ( .A(wk_share3[10]), .B(input3[10]), .Z(
        Midori_add_Result_Start3[10]) );
  XOR2_X1 Midori_U129 ( .A(wk_share3[0]), .B(input3[0]), .Z(
        Midori_add_Result_Start3[0]) );
  XOR2_X1 Midori_U128 ( .A(wk_share2[9]), .B(input2[9]), .Z(
        Midori_add_Result_Start2[9]) );
  XOR2_X1 Midori_U127 ( .A(wk_share2[8]), .B(input2[8]), .Z(
        Midori_add_Result_Start2[8]) );
  XOR2_X1 Midori_U126 ( .A(wk_share2[7]), .B(input2[7]), .Z(
        Midori_add_Result_Start2[7]) );
  XOR2_X1 Midori_U125 ( .A(wk_share2[6]), .B(input2[6]), .Z(
        Midori_add_Result_Start2[6]) );
  XOR2_X1 Midori_U124 ( .A(wk_share2[63]), .B(input2[63]), .Z(
        Midori_add_Result_Start2[63]) );
  XOR2_X1 Midori_U123 ( .A(wk_share2[62]), .B(input2[62]), .Z(
        Midori_add_Result_Start2[62]) );
  XOR2_X1 Midori_U122 ( .A(wk_share2[61]), .B(input2[61]), .Z(
        Midori_add_Result_Start2[61]) );
  XOR2_X1 Midori_U121 ( .A(wk_share2[60]), .B(input2[60]), .Z(
        Midori_add_Result_Start2[60]) );
  XOR2_X1 Midori_U120 ( .A(wk_share2[5]), .B(input2[5]), .Z(
        Midori_add_Result_Start2[5]) );
  XOR2_X1 Midori_U119 ( .A(wk_share2[59]), .B(input2[59]), .Z(
        Midori_add_Result_Start2[59]) );
  XOR2_X1 Midori_U118 ( .A(wk_share2[58]), .B(input2[58]), .Z(
        Midori_add_Result_Start2[58]) );
  XOR2_X1 Midori_U117 ( .A(wk_share2[57]), .B(input2[57]), .Z(
        Midori_add_Result_Start2[57]) );
  XOR2_X1 Midori_U116 ( .A(wk_share2[56]), .B(input2[56]), .Z(
        Midori_add_Result_Start2[56]) );
  XOR2_X1 Midori_U115 ( .A(wk_share2[55]), .B(input2[55]), .Z(
        Midori_add_Result_Start2[55]) );
  XOR2_X1 Midori_U114 ( .A(wk_share2[54]), .B(input2[54]), .Z(
        Midori_add_Result_Start2[54]) );
  XOR2_X1 Midori_U113 ( .A(wk_share2[53]), .B(input2[53]), .Z(
        Midori_add_Result_Start2[53]) );
  XOR2_X1 Midori_U112 ( .A(wk_share2[52]), .B(input2[52]), .Z(
        Midori_add_Result_Start2[52]) );
  XOR2_X1 Midori_U111 ( .A(wk_share2[51]), .B(input2[51]), .Z(
        Midori_add_Result_Start2[51]) );
  XOR2_X1 Midori_U110 ( .A(wk_share2[50]), .B(input2[50]), .Z(
        Midori_add_Result_Start2[50]) );
  XOR2_X1 Midori_U109 ( .A(wk_share2[4]), .B(input2[4]), .Z(
        Midori_add_Result_Start2[4]) );
  XOR2_X1 Midori_U108 ( .A(wk_share2[49]), .B(input2[49]), .Z(
        Midori_add_Result_Start2[49]) );
  XOR2_X1 Midori_U107 ( .A(wk_share2[48]), .B(input2[48]), .Z(
        Midori_add_Result_Start2[48]) );
  XOR2_X1 Midori_U106 ( .A(wk_share2[47]), .B(input2[47]), .Z(
        Midori_add_Result_Start2[47]) );
  XOR2_X1 Midori_U105 ( .A(wk_share2[46]), .B(input2[46]), .Z(
        Midori_add_Result_Start2[46]) );
  XOR2_X1 Midori_U104 ( .A(wk_share2[45]), .B(input2[45]), .Z(
        Midori_add_Result_Start2[45]) );
  XOR2_X1 Midori_U103 ( .A(wk_share2[44]), .B(input2[44]), .Z(
        Midori_add_Result_Start2[44]) );
  XOR2_X1 Midori_U102 ( .A(wk_share2[43]), .B(input2[43]), .Z(
        Midori_add_Result_Start2[43]) );
  XOR2_X1 Midori_U101 ( .A(wk_share2[42]), .B(input2[42]), .Z(
        Midori_add_Result_Start2[42]) );
  XOR2_X1 Midori_U100 ( .A(wk_share2[41]), .B(input2[41]), .Z(
        Midori_add_Result_Start2[41]) );
  XOR2_X1 Midori_U99 ( .A(wk_share2[40]), .B(input2[40]), .Z(
        Midori_add_Result_Start2[40]) );
  XOR2_X1 Midori_U98 ( .A(wk_share2[3]), .B(input2[3]), .Z(
        Midori_add_Result_Start2[3]) );
  XOR2_X1 Midori_U97 ( .A(wk_share2[39]), .B(input2[39]), .Z(
        Midori_add_Result_Start2[39]) );
  XOR2_X1 Midori_U96 ( .A(wk_share2[38]), .B(input2[38]), .Z(
        Midori_add_Result_Start2[38]) );
  XOR2_X1 Midori_U95 ( .A(wk_share2[37]), .B(input2[37]), .Z(
        Midori_add_Result_Start2[37]) );
  XOR2_X1 Midori_U94 ( .A(wk_share2[36]), .B(input2[36]), .Z(
        Midori_add_Result_Start2[36]) );
  XOR2_X1 Midori_U93 ( .A(wk_share2[35]), .B(input2[35]), .Z(
        Midori_add_Result_Start2[35]) );
  XOR2_X1 Midori_U92 ( .A(wk_share2[34]), .B(input2[34]), .Z(
        Midori_add_Result_Start2[34]) );
  XOR2_X1 Midori_U91 ( .A(wk_share2[33]), .B(input2[33]), .Z(
        Midori_add_Result_Start2[33]) );
  XOR2_X1 Midori_U90 ( .A(wk_share2[32]), .B(input2[32]), .Z(
        Midori_add_Result_Start2[32]) );
  XOR2_X1 Midori_U89 ( .A(wk_share2[31]), .B(input2[31]), .Z(
        Midori_add_Result_Start2[31]) );
  XOR2_X1 Midori_U88 ( .A(wk_share2[30]), .B(input2[30]), .Z(
        Midori_add_Result_Start2[30]) );
  XOR2_X1 Midori_U87 ( .A(wk_share2[2]), .B(input2[2]), .Z(
        Midori_add_Result_Start2[2]) );
  XOR2_X1 Midori_U86 ( .A(wk_share2[29]), .B(input2[29]), .Z(
        Midori_add_Result_Start2[29]) );
  XOR2_X1 Midori_U85 ( .A(wk_share2[28]), .B(input2[28]), .Z(
        Midori_add_Result_Start2[28]) );
  XOR2_X1 Midori_U84 ( .A(wk_share2[27]), .B(input2[27]), .Z(
        Midori_add_Result_Start2[27]) );
  XOR2_X1 Midori_U83 ( .A(wk_share2[26]), .B(input2[26]), .Z(
        Midori_add_Result_Start2[26]) );
  XOR2_X1 Midori_U82 ( .A(wk_share2[25]), .B(input2[25]), .Z(
        Midori_add_Result_Start2[25]) );
  XOR2_X1 Midori_U81 ( .A(wk_share2[24]), .B(input2[24]), .Z(
        Midori_add_Result_Start2[24]) );
  XOR2_X1 Midori_U80 ( .A(wk_share2[23]), .B(input2[23]), .Z(
        Midori_add_Result_Start2[23]) );
  XOR2_X1 Midori_U79 ( .A(wk_share2[22]), .B(input2[22]), .Z(
        Midori_add_Result_Start2[22]) );
  XOR2_X1 Midori_U78 ( .A(wk_share2[21]), .B(input2[21]), .Z(
        Midori_add_Result_Start2[21]) );
  XOR2_X1 Midori_U77 ( .A(wk_share2[20]), .B(input2[20]), .Z(
        Midori_add_Result_Start2[20]) );
  XOR2_X1 Midori_U76 ( .A(wk_share2[1]), .B(input2[1]), .Z(
        Midori_add_Result_Start2[1]) );
  XOR2_X1 Midori_U75 ( .A(wk_share2[19]), .B(input2[19]), .Z(
        Midori_add_Result_Start2[19]) );
  XOR2_X1 Midori_U74 ( .A(wk_share2[18]), .B(input2[18]), .Z(
        Midori_add_Result_Start2[18]) );
  XOR2_X1 Midori_U73 ( .A(wk_share2[17]), .B(input2[17]), .Z(
        Midori_add_Result_Start2[17]) );
  XOR2_X1 Midori_U72 ( .A(wk_share2[16]), .B(input2[16]), .Z(
        Midori_add_Result_Start2[16]) );
  XOR2_X1 Midori_U71 ( .A(wk_share2[15]), .B(input2[15]), .Z(
        Midori_add_Result_Start2[15]) );
  XOR2_X1 Midori_U70 ( .A(wk_share2[14]), .B(input2[14]), .Z(
        Midori_add_Result_Start2[14]) );
  XOR2_X1 Midori_U69 ( .A(wk_share2[13]), .B(input2[13]), .Z(
        Midori_add_Result_Start2[13]) );
  XOR2_X1 Midori_U68 ( .A(wk_share2[12]), .B(input2[12]), .Z(
        Midori_add_Result_Start2[12]) );
  XOR2_X1 Midori_U67 ( .A(wk_share2[11]), .B(input2[11]), .Z(
        Midori_add_Result_Start2[11]) );
  XOR2_X1 Midori_U66 ( .A(wk_share2[10]), .B(input2[10]), .Z(
        Midori_add_Result_Start2[10]) );
  XOR2_X1 Midori_U65 ( .A(wk_share2[0]), .B(input2[0]), .Z(
        Midori_add_Result_Start2[0]) );
  XOR2_X1 Midori_U64 ( .A(wk_share1[9]), .B(input1[9]), .Z(
        Midori_add_Result_Start1[9]) );
  XOR2_X1 Midori_U63 ( .A(wk_share1[8]), .B(input1[8]), .Z(
        Midori_add_Result_Start1[8]) );
  XOR2_X1 Midori_U62 ( .A(wk_share1[7]), .B(input1[7]), .Z(
        Midori_add_Result_Start1[7]) );
  XOR2_X1 Midori_U61 ( .A(wk_share1[6]), .B(input1[6]), .Z(
        Midori_add_Result_Start1[6]) );
  XOR2_X1 Midori_U60 ( .A(wk_share1[63]), .B(input1[63]), .Z(
        Midori_add_Result_Start1[63]) );
  XOR2_X1 Midori_U59 ( .A(wk_share1[62]), .B(input1[62]), .Z(
        Midori_add_Result_Start1[62]) );
  XOR2_X1 Midori_U58 ( .A(wk_share1[61]), .B(input1[61]), .Z(
        Midori_add_Result_Start1[61]) );
  XOR2_X1 Midori_U57 ( .A(wk_share1[60]), .B(input1[60]), .Z(
        Midori_add_Result_Start1[60]) );
  XOR2_X1 Midori_U56 ( .A(wk_share1[5]), .B(input1[5]), .Z(
        Midori_add_Result_Start1[5]) );
  XOR2_X1 Midori_U55 ( .A(wk_share1[59]), .B(input1[59]), .Z(
        Midori_add_Result_Start1[59]) );
  XOR2_X1 Midori_U54 ( .A(wk_share1[58]), .B(input1[58]), .Z(
        Midori_add_Result_Start1[58]) );
  XOR2_X1 Midori_U53 ( .A(wk_share1[57]), .B(input1[57]), .Z(
        Midori_add_Result_Start1[57]) );
  XOR2_X1 Midori_U52 ( .A(wk_share1[56]), .B(input1[56]), .Z(
        Midori_add_Result_Start1[56]) );
  XOR2_X1 Midori_U51 ( .A(wk_share1[55]), .B(input1[55]), .Z(
        Midori_add_Result_Start1[55]) );
  XOR2_X1 Midori_U50 ( .A(wk_share1[54]), .B(input1[54]), .Z(
        Midori_add_Result_Start1[54]) );
  XOR2_X1 Midori_U49 ( .A(wk_share1[53]), .B(input1[53]), .Z(
        Midori_add_Result_Start1[53]) );
  XOR2_X1 Midori_U48 ( .A(wk_share1[52]), .B(input1[52]), .Z(
        Midori_add_Result_Start1[52]) );
  XOR2_X1 Midori_U47 ( .A(wk_share1[51]), .B(input1[51]), .Z(
        Midori_add_Result_Start1[51]) );
  XOR2_X1 Midori_U46 ( .A(wk_share1[50]), .B(input1[50]), .Z(
        Midori_add_Result_Start1[50]) );
  XOR2_X1 Midori_U45 ( .A(wk_share1[4]), .B(input1[4]), .Z(
        Midori_add_Result_Start1[4]) );
  XOR2_X1 Midori_U44 ( .A(wk_share1[49]), .B(input1[49]), .Z(
        Midori_add_Result_Start1[49]) );
  XOR2_X1 Midori_U43 ( .A(wk_share1[48]), .B(input1[48]), .Z(
        Midori_add_Result_Start1[48]) );
  XOR2_X1 Midori_U42 ( .A(wk_share1[47]), .B(input1[47]), .Z(
        Midori_add_Result_Start1[47]) );
  XOR2_X1 Midori_U41 ( .A(wk_share1[46]), .B(input1[46]), .Z(
        Midori_add_Result_Start1[46]) );
  XOR2_X1 Midori_U40 ( .A(wk_share1[45]), .B(input1[45]), .Z(
        Midori_add_Result_Start1[45]) );
  XOR2_X1 Midori_U39 ( .A(wk_share1[44]), .B(input1[44]), .Z(
        Midori_add_Result_Start1[44]) );
  XOR2_X1 Midori_U38 ( .A(wk_share1[43]), .B(input1[43]), .Z(
        Midori_add_Result_Start1[43]) );
  XOR2_X1 Midori_U37 ( .A(wk_share1[42]), .B(input1[42]), .Z(
        Midori_add_Result_Start1[42]) );
  XOR2_X1 Midori_U36 ( .A(wk_share1[41]), .B(input1[41]), .Z(
        Midori_add_Result_Start1[41]) );
  XOR2_X1 Midori_U35 ( .A(wk_share1[40]), .B(input1[40]), .Z(
        Midori_add_Result_Start1[40]) );
  XOR2_X1 Midori_U34 ( .A(wk_share1[3]), .B(input1[3]), .Z(
        Midori_add_Result_Start1[3]) );
  XOR2_X1 Midori_U33 ( .A(wk_share1[39]), .B(input1[39]), .Z(
        Midori_add_Result_Start1[39]) );
  XOR2_X1 Midori_U32 ( .A(wk_share1[38]), .B(input1[38]), .Z(
        Midori_add_Result_Start1[38]) );
  XOR2_X1 Midori_U31 ( .A(wk_share1[37]), .B(input1[37]), .Z(
        Midori_add_Result_Start1[37]) );
  XOR2_X1 Midori_U30 ( .A(wk_share1[36]), .B(input1[36]), .Z(
        Midori_add_Result_Start1[36]) );
  XOR2_X1 Midori_U29 ( .A(wk_share1[35]), .B(input1[35]), .Z(
        Midori_add_Result_Start1[35]) );
  XOR2_X1 Midori_U28 ( .A(wk_share1[34]), .B(input1[34]), .Z(
        Midori_add_Result_Start1[34]) );
  XOR2_X1 Midori_U27 ( .A(wk_share1[33]), .B(input1[33]), .Z(
        Midori_add_Result_Start1[33]) );
  XOR2_X1 Midori_U26 ( .A(wk_share1[32]), .B(input1[32]), .Z(
        Midori_add_Result_Start1[32]) );
  XOR2_X1 Midori_U25 ( .A(wk_share1[31]), .B(input1[31]), .Z(
        Midori_add_Result_Start1[31]) );
  XOR2_X1 Midori_U24 ( .A(wk_share1[30]), .B(input1[30]), .Z(
        Midori_add_Result_Start1[30]) );
  XOR2_X1 Midori_U23 ( .A(wk_share1[2]), .B(input1[2]), .Z(
        Midori_add_Result_Start1[2]) );
  XOR2_X1 Midori_U22 ( .A(wk_share1[29]), .B(input1[29]), .Z(
        Midori_add_Result_Start1[29]) );
  XOR2_X1 Midori_U21 ( .A(wk_share1[28]), .B(input1[28]), .Z(
        Midori_add_Result_Start1[28]) );
  XOR2_X1 Midori_U20 ( .A(wk_share1[27]), .B(input1[27]), .Z(
        Midori_add_Result_Start1[27]) );
  XOR2_X1 Midori_U19 ( .A(wk_share1[26]), .B(input1[26]), .Z(
        Midori_add_Result_Start1[26]) );
  XOR2_X1 Midori_U18 ( .A(wk_share1[25]), .B(input1[25]), .Z(
        Midori_add_Result_Start1[25]) );
  XOR2_X1 Midori_U17 ( .A(wk_share1[24]), .B(input1[24]), .Z(
        Midori_add_Result_Start1[24]) );
  XOR2_X1 Midori_U16 ( .A(wk_share1[23]), .B(input1[23]), .Z(
        Midori_add_Result_Start1[23]) );
  XOR2_X1 Midori_U15 ( .A(wk_share1[22]), .B(input1[22]), .Z(
        Midori_add_Result_Start1[22]) );
  XOR2_X1 Midori_U14 ( .A(wk_share1[21]), .B(input1[21]), .Z(
        Midori_add_Result_Start1[21]) );
  XOR2_X1 Midori_U13 ( .A(wk_share1[20]), .B(input1[20]), .Z(
        Midori_add_Result_Start1[20]) );
  XOR2_X1 Midori_U12 ( .A(wk_share1[1]), .B(input1[1]), .Z(
        Midori_add_Result_Start1[1]) );
  XOR2_X1 Midori_U11 ( .A(wk_share1[19]), .B(input1[19]), .Z(
        Midori_add_Result_Start1[19]) );
  XOR2_X1 Midori_U10 ( .A(wk_share1[18]), .B(input1[18]), .Z(
        Midori_add_Result_Start1[18]) );
  XOR2_X1 Midori_U9 ( .A(wk_share1[17]), .B(input1[17]), .Z(
        Midori_add_Result_Start1[17]) );
  XOR2_X1 Midori_U8 ( .A(wk_share1[16]), .B(input1[16]), .Z(
        Midori_add_Result_Start1[16]) );
  XOR2_X1 Midori_U7 ( .A(wk_share1[15]), .B(input1[15]), .Z(
        Midori_add_Result_Start1[15]) );
  XOR2_X1 Midori_U6 ( .A(wk_share1[14]), .B(input1[14]), .Z(
        Midori_add_Result_Start1[14]) );
  XOR2_X1 Midori_U5 ( .A(wk_share1[13]), .B(input1[13]), .Z(
        Midori_add_Result_Start1[13]) );
  XOR2_X1 Midori_U4 ( .A(wk_share1[12]), .B(input1[12]), .Z(
        Midori_add_Result_Start1[12]) );
  XOR2_X1 Midori_U3 ( .A(wk_share1[11]), .B(input1[11]), .Z(
        Midori_add_Result_Start1[11]) );
  XOR2_X1 Midori_U2 ( .A(wk_share1[10]), .B(input1[10]), .Z(
        Midori_add_Result_Start1[10]) );
  XOR2_X1 Midori_U1 ( .A(wk_share1[0]), .B(input1[0]), .Z(
        Midori_add_Result_Start1[0]) );
  OAI21_X1 Midori_rounds_U1213 ( .B1(Midori_rounds_n2067), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2065), .ZN(
        Midori_rounds_sub_Sub_0_S1_InAff_out1[1]) );
  AOI22_X1 Midori_rounds_U1212 ( .A1(reset), .A2(Midori_add_Result_Start1[0]), 
        .B1(Midori_rounds_n2064), .B2(Midori_rounds_SR_Inv_Result1[0]), .ZN(
        Midori_rounds_n2065) );
  XOR2_X1 Midori_rounds_U1211 ( .A(Midori_rounds_SR_Inv_Result1[28]), .B(
        Midori_rounds_n2063), .Z(Midori_rounds_n2067) );
  OAI21_X1 Midori_rounds_U1210 ( .B1(Midori_rounds_n2062), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2061), .ZN(
        Midori_rounds_sub_Sub_0_S2_InAff_out1[1]) );
  AOI22_X1 Midori_rounds_U1209 ( .A1(reset), .A2(Midori_add_Result_Start1[4]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result1[4]), .ZN(
        Midori_rounds_n2061) );
  XOR2_X1 Midori_rounds_U1208 ( .A(Midori_rounds_SR_Inv_Result1[52]), .B(
        Midori_rounds_n2060), .Z(Midori_rounds_n2062) );
  OAI21_X1 Midori_rounds_U1207 ( .B1(Midori_rounds_n2059), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2058), .ZN(
        Midori_rounds_sub_Sub_1_S1_InAff_out1[1]) );
  AOI22_X1 Midori_rounds_U1206 ( .A1(reset), .A2(Midori_add_Result_Start1[8]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result1[8]), .ZN(
        Midori_rounds_n2058) );
  XOR2_X1 Midori_rounds_U1205 ( .A(Midori_rounds_SR_Inv_Result1[8]), .B(
        Midori_rounds_n2057), .Z(Midori_rounds_n2059) );
  OAI21_X1 Midori_rounds_U1204 ( .B1(Midori_rounds_n2056), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2055), .ZN(
        Midori_rounds_sub_Sub_1_S2_InAff_out1[1]) );
  AOI22_X1 Midori_rounds_U1203 ( .A1(reset), .A2(Midori_add_Result_Start1[12]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[12]), .ZN(
        Midori_rounds_n2055) );
  XOR2_X1 Midori_rounds_U1202 ( .A(Midori_rounds_SR_Inv_Result1[32]), .B(
        Midori_rounds_n2054), .Z(Midori_rounds_n2056) );
  OAI21_X1 Midori_rounds_U1201 ( .B1(Midori_rounds_n2053), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2052), .ZN(
        Midori_rounds_sub_Sub_2_S1_InAff_out1[1]) );
  AOI22_X1 Midori_rounds_U1200 ( .A1(reset), .A2(Midori_add_Result_Start1[16]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result1[16]), .ZN(
        Midori_rounds_n2052) );
  XOR2_X1 Midori_rounds_U1199 ( .A(Midori_rounds_SR_Inv_Result1[36]), .B(
        Midori_rounds_n2051), .Z(Midori_rounds_n2053) );
  OAI21_X1 Midori_rounds_U1198 ( .B1(Midori_rounds_n2050), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2049), .ZN(
        Midori_rounds_sub_Sub_2_S2_InAff_out1[1]) );
  AOI22_X1 Midori_rounds_U1197 ( .A1(reset), .A2(Midori_add_Result_Start1[20]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result1[20]), .ZN(
        Midori_rounds_n2049) );
  XOR2_X1 Midori_rounds_U1196 ( .A(Midori_rounds_SR_Inv_Result1[12]), .B(
        Midori_rounds_n2048), .Z(Midori_rounds_n2050) );
  OAI21_X1 Midori_rounds_U1195 ( .B1(Midori_rounds_n2047), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2046), .ZN(
        Midori_rounds_sub_Sub_3_S1_InAff_out1[1]) );
  AOI22_X1 Midori_rounds_U1194 ( .A1(reset), .A2(Midori_add_Result_Start1[24]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result1[24]), .ZN(
        Midori_rounds_n2046) );
  XOR2_X1 Midori_rounds_U1193 ( .A(Midori_rounds_SR_Inv_Result1[48]), .B(
        Midori_rounds_n2045), .Z(Midori_rounds_n2047) );
  OAI21_X1 Midori_rounds_U1192 ( .B1(Midori_rounds_n2044), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2043), .ZN(
        Midori_rounds_sub_Sub_3_S2_InAff_out1[1]) );
  AOI22_X1 Midori_rounds_U1191 ( .A1(reset), .A2(Midori_add_Result_Start1[28]), 
        .B1(Midori_rounds_n2064), .B2(Midori_rounds_SR_Inv_Result1[28]), .ZN(
        Midori_rounds_n2043) );
  XOR2_X1 Midori_rounds_U1190 ( .A(Midori_rounds_SR_Inv_Result1[24]), .B(
        Midori_rounds_n2042), .Z(Midori_rounds_n2044) );
  OAI21_X1 Midori_rounds_U1189 ( .B1(Midori_rounds_n2041), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2040), .ZN(
        Midori_rounds_sub_Sub_4_S1_InAff_out1[1]) );
  AOI22_X1 Midori_rounds_U1188 ( .A1(reset), .A2(Midori_add_Result_Start1[32]), 
        .B1(Midori_rounds_n2064), .B2(Midori_rounds_SR_Inv_Result1[32]), .ZN(
        Midori_rounds_n2040) );
  XOR2_X1 Midori_rounds_U1187 ( .A(Midori_rounds_SR_Inv_Result1[56]), .B(
        Midori_rounds_n2039), .Z(Midori_rounds_n2041) );
  OAI21_X1 Midori_rounds_U1186 ( .B1(Midori_rounds_n2038), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2037), .ZN(
        Midori_rounds_sub_Sub_4_S2_InAff_out1[1]) );
  AOI22_X1 Midori_rounds_U1185 ( .A1(reset), .A2(Midori_add_Result_Start1[36]), 
        .B1(Midori_rounds_n2064), .B2(Midori_rounds_SR_Inv_Result1[36]), .ZN(
        Midori_rounds_n2037) );
  XOR2_X1 Midori_rounds_U1184 ( .A(Midori_rounds_SR_Inv_Result1[16]), .B(
        Midori_rounds_n2036), .Z(Midori_rounds_n2038) );
  OAI21_X1 Midori_rounds_U1183 ( .B1(Midori_rounds_n2035), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2034), .ZN(
        Midori_rounds_sub_Sub_5_S1_InAff_out1[1]) );
  AOI22_X1 Midori_rounds_U1182 ( .A1(reset), .A2(Midori_add_Result_Start1[40]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result1[40]), .ZN(
        Midori_rounds_n2034) );
  XOR2_X1 Midori_rounds_U1181 ( .A(Midori_rounds_SR_Inv_Result1[44]), .B(
        Midori_rounds_n2033), .Z(Midori_rounds_n2035) );
  OAI21_X1 Midori_rounds_U1180 ( .B1(Midori_rounds_n2032), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n2031), .ZN(
        Midori_rounds_sub_Sub_5_S2_InAff_out1[1]) );
  AOI22_X1 Midori_rounds_U1179 ( .A1(reset), .A2(Midori_add_Result_Start1[44]), 
        .B1(Midori_rounds_n2064), .B2(Midori_rounds_SR_Inv_Result1[44]), .ZN(
        Midori_rounds_n2031) );
  XOR2_X1 Midori_rounds_U1178 ( .A(Midori_rounds_SR_Inv_Result1[4]), .B(
        Midori_rounds_n2030), .Z(Midori_rounds_n2032) );
  OAI21_X1 Midori_rounds_U1177 ( .B1(Midori_rounds_n2029), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2028), .ZN(
        Midori_rounds_sub_Sub_6_S1_InAff_out1[1]) );
  AOI22_X1 Midori_rounds_U1176 ( .A1(reset), .A2(Midori_add_Result_Start1[48]), 
        .B1(Midori_rounds_n2064), .B2(Midori_rounds_SR_Inv_Result1[48]), .ZN(
        Midori_rounds_n2028) );
  XOR2_X1 Midori_rounds_U1175 ( .A(Midori_rounds_SR_Inv_Result1[0]), .B(
        Midori_rounds_n2027), .Z(Midori_rounds_n2029) );
  OAI21_X1 Midori_rounds_U1174 ( .B1(Midori_rounds_n2026), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2025), .ZN(
        Midori_rounds_sub_Sub_6_S2_InAff_out1[1]) );
  AOI22_X1 Midori_rounds_U1173 ( .A1(reset), .A2(Midori_add_Result_Start1[52]), 
        .B1(Midori_rounds_n2064), .B2(Midori_rounds_SR_Inv_Result1[52]), .ZN(
        Midori_rounds_n2025) );
  XOR2_X1 Midori_rounds_U1172 ( .A(Midori_rounds_SR_Inv_Result1[40]), .B(
        Midori_rounds_n2024), .Z(Midori_rounds_n2026) );
  OAI21_X1 Midori_rounds_U1171 ( .B1(Midori_rounds_n2023), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2022), .ZN(
        Midori_rounds_sub_Sub_7_S1_InAff_out1[1]) );
  AOI22_X1 Midori_rounds_U1170 ( .A1(reset), .A2(Midori_add_Result_Start1[56]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result1[56]), .ZN(
        Midori_rounds_n2022) );
  XOR2_X1 Midori_rounds_U1169 ( .A(Midori_rounds_SR_Inv_Result1[20]), .B(
        Midori_rounds_n2021), .Z(Midori_rounds_n2023) );
  OAI21_X1 Midori_rounds_U1168 ( .B1(Midori_rounds_n2020), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2019), .ZN(
        Midori_rounds_sub_Sub_7_S2_InAff_out1[1]) );
  AOI22_X1 Midori_rounds_U1167 ( .A1(reset), .A2(Midori_add_Result_Start1[60]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result1[60]), .ZN(
        Midori_rounds_n2019) );
  XOR2_X1 Midori_rounds_U1166 ( .A(Midori_rounds_SR_Inv_Result1[60]), .B(
        Midori_rounds_n2018), .Z(Midori_rounds_n2020) );
  OAI21_X1 Midori_rounds_U1165 ( .B1(Midori_rounds_n2017), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2016), .ZN(
        Midori_rounds_sub_Sub_0_S1_InAff_out1[0]) );
  AOI22_X1 Midori_rounds_U1164 ( .A1(reset), .A2(Midori_add_Result_Start1[1]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result1[1]), .ZN(
        Midori_rounds_n2016) );
  XOR2_X1 Midori_rounds_U1163 ( .A(Midori_rounds_SR_Inv_Result1[29]), .B(
        Midori_rounds_n2015), .Z(Midori_rounds_n2017) );
  OAI21_X1 Midori_rounds_U1162 ( .B1(Midori_rounds_n2014), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2013), .ZN(Midori_rounds_n806)
         );
  AOI22_X1 Midori_rounds_U1161 ( .A1(reset), .A2(Midori_add_Result_Start1[2]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result1[2]), .ZN(
        Midori_rounds_n2013) );
  XOR2_X1 Midori_rounds_U1160 ( .A(Midori_rounds_SR_Inv_Result1[30]), .B(
        Midori_rounds_n2012), .Z(Midori_rounds_n2014) );
  OAI21_X1 Midori_rounds_U1159 ( .B1(Midori_rounds_n2011), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2010), .ZN(
        Midori_rounds_sub_Sub_0_S1_InAff_out1[2]) );
  AOI22_X1 Midori_rounds_U1158 ( .A1(reset), .A2(Midori_add_Result_Start1[3]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result1[3]), .ZN(
        Midori_rounds_n2010) );
  XOR2_X1 Midori_rounds_U1157 ( .A(Midori_rounds_SR_Inv_Result1[31]), .B(
        Midori_rounds_n2009), .Z(Midori_rounds_n2011) );
  OAI21_X1 Midori_rounds_U1156 ( .B1(Midori_rounds_n2008), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2007), .ZN(
        Midori_rounds_sub_Sub_0_S2_InAff_out1[0]) );
  AOI22_X1 Midori_rounds_U1155 ( .A1(reset), .A2(Midori_add_Result_Start1[5]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result1[5]), .ZN(
        Midori_rounds_n2007) );
  XOR2_X1 Midori_rounds_U1154 ( .A(Midori_rounds_SR_Inv_Result1[53]), .B(
        Midori_rounds_n2006), .Z(Midori_rounds_n2008) );
  OAI21_X1 Midori_rounds_U1153 ( .B1(Midori_rounds_n2005), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2004), .ZN(Midori_rounds_n809)
         );
  AOI22_X1 Midori_rounds_U1152 ( .A1(reset), .A2(Midori_add_Result_Start1[6]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[6]), .ZN(
        Midori_rounds_n2004) );
  XOR2_X1 Midori_rounds_U1151 ( .A(Midori_rounds_SR_Inv_Result1[54]), .B(
        Midori_rounds_n2003), .Z(Midori_rounds_n2005) );
  OAI21_X1 Midori_rounds_U1150 ( .B1(Midori_rounds_n2002), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n2001), .ZN(
        Midori_rounds_sub_Sub_0_S2_InAff_out1[2]) );
  AOI22_X1 Midori_rounds_U1149 ( .A1(reset), .A2(Midori_add_Result_Start1[7]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result1[7]), .ZN(
        Midori_rounds_n2001) );
  XOR2_X1 Midori_rounds_U1148 ( .A(Midori_rounds_SR_Inv_Result1[55]), .B(
        Midori_rounds_n2000), .Z(Midori_rounds_n2002) );
  OAI21_X1 Midori_rounds_U1147 ( .B1(Midori_rounds_n1999), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1998), .ZN(
        Midori_rounds_sub_Sub_1_S1_InAff_out1[0]) );
  AOI22_X1 Midori_rounds_U1146 ( .A1(reset), .A2(Midori_add_Result_Start1[9]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result1[9]), .ZN(
        Midori_rounds_n1998) );
  XOR2_X1 Midori_rounds_U1145 ( .A(Midori_rounds_SR_Inv_Result1[9]), .B(
        Midori_rounds_n1997), .Z(Midori_rounds_n1999) );
  OAI21_X1 Midori_rounds_U1144 ( .B1(Midori_rounds_n1996), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1995), .ZN(Midori_rounds_n812)
         );
  AOI22_X1 Midori_rounds_U1143 ( .A1(reset), .A2(Midori_add_Result_Start1[10]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result1[10]), .ZN(
        Midori_rounds_n1995) );
  XOR2_X1 Midori_rounds_U1142 ( .A(Midori_rounds_SR_Inv_Result1[10]), .B(
        Midori_rounds_n1994), .Z(Midori_rounds_n1996) );
  OAI21_X1 Midori_rounds_U1141 ( .B1(Midori_rounds_n1993), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1992), .ZN(
        Midori_rounds_sub_Sub_1_S1_InAff_out1[2]) );
  AOI22_X1 Midori_rounds_U1140 ( .A1(reset), .A2(Midori_add_Result_Start1[11]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[11]), .ZN(
        Midori_rounds_n1992) );
  XOR2_X1 Midori_rounds_U1139 ( .A(Midori_rounds_SR_Inv_Result1[11]), .B(
        Midori_rounds_n1991), .Z(Midori_rounds_n1993) );
  OAI21_X1 Midori_rounds_U1138 ( .B1(Midori_rounds_n1990), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1989), .ZN(
        Midori_rounds_sub_Sub_1_S2_InAff_out1[0]) );
  AOI22_X1 Midori_rounds_U1137 ( .A1(reset), .A2(Midori_add_Result_Start1[13]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[13]), .ZN(
        Midori_rounds_n1989) );
  XOR2_X1 Midori_rounds_U1136 ( .A(Midori_rounds_SR_Inv_Result1[33]), .B(
        Midori_rounds_n1988), .Z(Midori_rounds_n1990) );
  OAI21_X1 Midori_rounds_U1135 ( .B1(Midori_rounds_n1987), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1986), .ZN(Midori_rounds_n815)
         );
  AOI22_X1 Midori_rounds_U1134 ( .A1(reset), .A2(Midori_add_Result_Start1[14]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[14]), .ZN(
        Midori_rounds_n1986) );
  XOR2_X1 Midori_rounds_U1133 ( .A(Midori_rounds_SR_Inv_Result1[34]), .B(
        Midori_rounds_n1985), .Z(Midori_rounds_n1987) );
  OAI21_X1 Midori_rounds_U1132 ( .B1(Midori_rounds_n1984), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1983), .ZN(
        Midori_rounds_sub_Sub_1_S2_InAff_out1[2]) );
  AOI22_X1 Midori_rounds_U1131 ( .A1(reset), .A2(Midori_add_Result_Start1[15]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[15]), .ZN(
        Midori_rounds_n1983) );
  XOR2_X1 Midori_rounds_U1130 ( .A(Midori_rounds_SR_Inv_Result1[35]), .B(
        Midori_rounds_n1982), .Z(Midori_rounds_n1984) );
  OAI21_X1 Midori_rounds_U1129 ( .B1(Midori_rounds_n1981), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1980), .ZN(
        Midori_rounds_sub_Sub_2_S1_InAff_out1[0]) );
  AOI22_X1 Midori_rounds_U1128 ( .A1(reset), .A2(Midori_add_Result_Start1[17]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[17]), .ZN(
        Midori_rounds_n1980) );
  XOR2_X1 Midori_rounds_U1127 ( .A(Midori_rounds_SR_Inv_Result1[37]), .B(
        Midori_rounds_n1979), .Z(Midori_rounds_n1981) );
  OAI21_X1 Midori_rounds_U1126 ( .B1(Midori_rounds_n1978), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1977), .ZN(Midori_rounds_n818)
         );
  AOI22_X1 Midori_rounds_U1125 ( .A1(reset), .A2(Midori_add_Result_Start1[18]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[18]), .ZN(
        Midori_rounds_n1977) );
  XOR2_X1 Midori_rounds_U1124 ( .A(Midori_rounds_SR_Inv_Result1[38]), .B(
        Midori_rounds_n1976), .Z(Midori_rounds_n1978) );
  OAI21_X1 Midori_rounds_U1123 ( .B1(Midori_rounds_n1975), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1974), .ZN(
        Midori_rounds_sub_Sub_2_S1_InAff_out1[2]) );
  AOI22_X1 Midori_rounds_U1122 ( .A1(reset), .A2(Midori_add_Result_Start1[19]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[19]), .ZN(
        Midori_rounds_n1974) );
  XOR2_X1 Midori_rounds_U1121 ( .A(Midori_rounds_SR_Inv_Result1[39]), .B(
        Midori_rounds_n1973), .Z(Midori_rounds_n1975) );
  OAI21_X1 Midori_rounds_U1120 ( .B1(Midori_rounds_n1972), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1971), .ZN(
        Midori_rounds_sub_Sub_2_S2_InAff_out1[0]) );
  AOI22_X1 Midori_rounds_U1119 ( .A1(reset), .A2(Midori_add_Result_Start1[21]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[21]), .ZN(
        Midori_rounds_n1971) );
  XOR2_X1 Midori_rounds_U1118 ( .A(Midori_rounds_SR_Inv_Result1[13]), .B(
        Midori_rounds_n1970), .Z(Midori_rounds_n1972) );
  OAI21_X1 Midori_rounds_U1117 ( .B1(Midori_rounds_n1969), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1968), .ZN(Midori_rounds_n821)
         );
  AOI22_X1 Midori_rounds_U1116 ( .A1(reset), .A2(Midori_add_Result_Start1[22]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[22]), .ZN(
        Midori_rounds_n1968) );
  XOR2_X1 Midori_rounds_U1115 ( .A(Midori_rounds_SR_Inv_Result1[14]), .B(
        Midori_rounds_n1967), .Z(Midori_rounds_n1969) );
  OAI21_X1 Midori_rounds_U1114 ( .B1(Midori_rounds_n1966), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1965), .ZN(
        Midori_rounds_sub_Sub_2_S2_InAff_out1[2]) );
  AOI22_X1 Midori_rounds_U1113 ( .A1(reset), .A2(Midori_add_Result_Start1[23]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[23]), .ZN(
        Midori_rounds_n1965) );
  XOR2_X1 Midori_rounds_U1112 ( .A(Midori_rounds_SR_Inv_Result1[15]), .B(
        Midori_rounds_n1964), .Z(Midori_rounds_n1966) );
  OAI21_X1 Midori_rounds_U1111 ( .B1(Midori_rounds_n1963), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1962), .ZN(
        Midori_rounds_sub_Sub_3_S1_InAff_out1[0]) );
  AOI22_X1 Midori_rounds_U1110 ( .A1(reset), .A2(Midori_add_Result_Start1[25]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[25]), .ZN(
        Midori_rounds_n1962) );
  XOR2_X1 Midori_rounds_U1109 ( .A(Midori_rounds_SR_Inv_Result1[49]), .B(
        Midori_rounds_n1961), .Z(Midori_rounds_n1963) );
  OAI21_X1 Midori_rounds_U1108 ( .B1(Midori_rounds_n1960), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1959), .ZN(Midori_rounds_n824)
         );
  AOI22_X1 Midori_rounds_U1107 ( .A1(reset), .A2(Midori_add_Result_Start1[26]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[26]), .ZN(
        Midori_rounds_n1959) );
  XOR2_X1 Midori_rounds_U1106 ( .A(Midori_rounds_SR_Inv_Result1[50]), .B(
        Midori_rounds_n1958), .Z(Midori_rounds_n1960) );
  OAI21_X1 Midori_rounds_U1105 ( .B1(Midori_rounds_n1957), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1956), .ZN(
        Midori_rounds_sub_Sub_3_S1_InAff_out1[2]) );
  AOI22_X1 Midori_rounds_U1104 ( .A1(reset), .A2(Midori_add_Result_Start1[27]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result1[27]), .ZN(
        Midori_rounds_n1956) );
  XOR2_X1 Midori_rounds_U1103 ( .A(Midori_rounds_SR_Inv_Result1[51]), .B(
        Midori_rounds_n1955), .Z(Midori_rounds_n1957) );
  OAI21_X1 Midori_rounds_U1102 ( .B1(Midori_rounds_n1954), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1953), .ZN(
        Midori_rounds_sub_Sub_3_S2_InAff_out1[0]) );
  AOI22_X1 Midori_rounds_U1101 ( .A1(reset), .A2(Midori_add_Result_Start1[29]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result1[29]), .ZN(
        Midori_rounds_n1953) );
  XOR2_X1 Midori_rounds_U1100 ( .A(Midori_rounds_SR_Inv_Result1[25]), .B(
        Midori_rounds_n1952), .Z(Midori_rounds_n1954) );
  OAI21_X1 Midori_rounds_U1099 ( .B1(Midori_rounds_n1951), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1950), .ZN(Midori_rounds_n827)
         );
  AOI22_X1 Midori_rounds_U1098 ( .A1(reset), .A2(Midori_add_Result_Start1[30]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result1[30]), .ZN(
        Midori_rounds_n1950) );
  XOR2_X1 Midori_rounds_U1097 ( .A(Midori_rounds_SR_Inv_Result1[26]), .B(
        Midori_rounds_n1949), .Z(Midori_rounds_n1951) );
  OAI21_X1 Midori_rounds_U1096 ( .B1(Midori_rounds_n1948), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1947), .ZN(
        Midori_rounds_sub_Sub_3_S2_InAff_out1[2]) );
  AOI22_X1 Midori_rounds_U1095 ( .A1(reset), .A2(Midori_add_Result_Start1[31]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result1[31]), .ZN(
        Midori_rounds_n1947) );
  XOR2_X1 Midori_rounds_U1094 ( .A(Midori_rounds_SR_Inv_Result1[27]), .B(
        Midori_rounds_n1946), .Z(Midori_rounds_n1948) );
  OAI21_X1 Midori_rounds_U1093 ( .B1(Midori_rounds_n1945), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1944), .ZN(
        Midori_rounds_sub_Sub_4_S1_InAff_out1[0]) );
  AOI22_X1 Midori_rounds_U1092 ( .A1(reset), .A2(Midori_add_Result_Start1[33]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result1[33]), .ZN(
        Midori_rounds_n1944) );
  XOR2_X1 Midori_rounds_U1091 ( .A(Midori_rounds_SR_Inv_Result1[57]), .B(
        Midori_rounds_n1943), .Z(Midori_rounds_n1945) );
  OAI21_X1 Midori_rounds_U1090 ( .B1(Midori_rounds_n1942), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1941), .ZN(Midori_rounds_n830)
         );
  AOI22_X1 Midori_rounds_U1089 ( .A1(reset), .A2(Midori_add_Result_Start1[34]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result1[34]), .ZN(
        Midori_rounds_n1941) );
  XOR2_X1 Midori_rounds_U1088 ( .A(Midori_rounds_SR_Inv_Result1[58]), .B(
        Midori_rounds_n1940), .Z(Midori_rounds_n1942) );
  OAI21_X1 Midori_rounds_U1087 ( .B1(Midori_rounds_n1939), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1938), .ZN(
        Midori_rounds_sub_Sub_4_S1_InAff_out1[2]) );
  AOI22_X1 Midori_rounds_U1086 ( .A1(reset), .A2(Midori_add_Result_Start1[35]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result1[35]), .ZN(
        Midori_rounds_n1938) );
  XOR2_X1 Midori_rounds_U1085 ( .A(Midori_rounds_SR_Inv_Result1[59]), .B(
        Midori_rounds_n1937), .Z(Midori_rounds_n1939) );
  OAI21_X1 Midori_rounds_U1084 ( .B1(Midori_rounds_n1936), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1935), .ZN(
        Midori_rounds_sub_Sub_4_S2_InAff_out1[0]) );
  AOI22_X1 Midori_rounds_U1083 ( .A1(reset), .A2(Midori_add_Result_Start1[37]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result1[37]), .ZN(
        Midori_rounds_n1935) );
  XOR2_X1 Midori_rounds_U1082 ( .A(Midori_rounds_SR_Inv_Result1[17]), .B(
        Midori_rounds_n1934), .Z(Midori_rounds_n1936) );
  OAI21_X1 Midori_rounds_U1081 ( .B1(Midori_rounds_n1933), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1932), .ZN(Midori_rounds_n833)
         );
  AOI22_X1 Midori_rounds_U1080 ( .A1(reset), .A2(Midori_add_Result_Start1[38]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[38]), .ZN(
        Midori_rounds_n1932) );
  XOR2_X1 Midori_rounds_U1079 ( .A(Midori_rounds_SR_Inv_Result1[18]), .B(
        Midori_rounds_n1931), .Z(Midori_rounds_n1933) );
  OAI21_X1 Midori_rounds_U1078 ( .B1(Midori_rounds_n1930), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1929), .ZN(
        Midori_rounds_sub_Sub_4_S2_InAff_out1[2]) );
  AOI22_X1 Midori_rounds_U1077 ( .A1(reset), .A2(Midori_add_Result_Start1[39]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result1[39]), .ZN(
        Midori_rounds_n1929) );
  XOR2_X1 Midori_rounds_U1076 ( .A(Midori_rounds_SR_Inv_Result1[19]), .B(
        Midori_rounds_n1928), .Z(Midori_rounds_n1930) );
  OAI21_X1 Midori_rounds_U1075 ( .B1(Midori_rounds_n1927), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1926), .ZN(
        Midori_rounds_sub_Sub_5_S1_InAff_out1[0]) );
  AOI22_X1 Midori_rounds_U1074 ( .A1(reset), .A2(Midori_add_Result_Start1[41]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result1[41]), .ZN(
        Midori_rounds_n1926) );
  XOR2_X1 Midori_rounds_U1073 ( .A(Midori_rounds_SR_Inv_Result1[45]), .B(
        Midori_rounds_n1925), .Z(Midori_rounds_n1927) );
  OAI21_X1 Midori_rounds_U1072 ( .B1(Midori_rounds_n1924), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1923), .ZN(Midori_rounds_n836)
         );
  AOI22_X1 Midori_rounds_U1071 ( .A1(reset), .A2(Midori_add_Result_Start1[42]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result1[42]), .ZN(
        Midori_rounds_n1923) );
  XOR2_X1 Midori_rounds_U1070 ( .A(Midori_rounds_SR_Inv_Result1[46]), .B(
        Midori_rounds_n1922), .Z(Midori_rounds_n1924) );
  OAI21_X1 Midori_rounds_U1069 ( .B1(Midori_rounds_n1921), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1920), .ZN(
        Midori_rounds_sub_Sub_5_S1_InAff_out1[2]) );
  AOI22_X1 Midori_rounds_U1068 ( .A1(reset), .A2(Midori_add_Result_Start1[43]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result1[43]), .ZN(
        Midori_rounds_n1920) );
  XOR2_X1 Midori_rounds_U1067 ( .A(Midori_rounds_SR_Inv_Result1[47]), .B(
        Midori_rounds_n1919), .Z(Midori_rounds_n1921) );
  OAI21_X1 Midori_rounds_U1066 ( .B1(Midori_rounds_n1918), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1917), .ZN(
        Midori_rounds_sub_Sub_5_S2_InAff_out1[0]) );
  AOI22_X1 Midori_rounds_U1065 ( .A1(reset), .A2(Midori_add_Result_Start1[45]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result1[45]), .ZN(
        Midori_rounds_n1917) );
  XOR2_X1 Midori_rounds_U1064 ( .A(Midori_rounds_SR_Inv_Result1[5]), .B(
        Midori_rounds_n1916), .Z(Midori_rounds_n1918) );
  OAI21_X1 Midori_rounds_U1063 ( .B1(Midori_rounds_n1915), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1914), .ZN(Midori_rounds_n839)
         );
  AOI22_X1 Midori_rounds_U1062 ( .A1(reset), .A2(Midori_add_Result_Start1[46]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result1[46]), .ZN(
        Midori_rounds_n1914) );
  XOR2_X1 Midori_rounds_U1061 ( .A(Midori_rounds_SR_Inv_Result1[6]), .B(
        Midori_rounds_n1913), .Z(Midori_rounds_n1915) );
  OAI21_X1 Midori_rounds_U1060 ( .B1(Midori_rounds_n1912), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1911), .ZN(
        Midori_rounds_sub_Sub_5_S2_InAff_out1[2]) );
  AOI22_X1 Midori_rounds_U1059 ( .A1(reset), .A2(Midori_add_Result_Start1[47]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result1[47]), .ZN(
        Midori_rounds_n1911) );
  XOR2_X1 Midori_rounds_U1058 ( .A(Midori_rounds_SR_Inv_Result1[7]), .B(
        Midori_rounds_n1910), .Z(Midori_rounds_n1912) );
  OAI21_X1 Midori_rounds_U1057 ( .B1(Midori_rounds_n1909), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1908), .ZN(
        Midori_rounds_sub_Sub_6_S1_InAff_out1[0]) );
  AOI22_X1 Midori_rounds_U1056 ( .A1(reset), .A2(Midori_add_Result_Start1[49]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result1[49]), .ZN(
        Midori_rounds_n1908) );
  XOR2_X1 Midori_rounds_U1055 ( .A(Midori_rounds_SR_Inv_Result1[1]), .B(
        Midori_rounds_n1907), .Z(Midori_rounds_n1909) );
  OAI21_X1 Midori_rounds_U1054 ( .B1(Midori_rounds_n1906), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1905), .ZN(Midori_rounds_n842)
         );
  AOI22_X1 Midori_rounds_U1053 ( .A1(reset), .A2(Midori_add_Result_Start1[50]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result1[50]), .ZN(
        Midori_rounds_n1905) );
  XOR2_X1 Midori_rounds_U1052 ( .A(Midori_rounds_SR_Inv_Result1[2]), .B(
        Midori_rounds_n1904), .Z(Midori_rounds_n1906) );
  OAI21_X1 Midori_rounds_U1051 ( .B1(Midori_rounds_n1903), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1902), .ZN(
        Midori_rounds_sub_Sub_6_S1_InAff_out1[2]) );
  AOI22_X1 Midori_rounds_U1050 ( .A1(reset), .A2(Midori_add_Result_Start1[51]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result1[51]), .ZN(
        Midori_rounds_n1902) );
  XOR2_X1 Midori_rounds_U1049 ( .A(Midori_rounds_SR_Inv_Result1[3]), .B(
        Midori_rounds_n1901), .Z(Midori_rounds_n1903) );
  OAI21_X1 Midori_rounds_U1048 ( .B1(Midori_rounds_n1900), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1899), .ZN(
        Midori_rounds_sub_Sub_6_S2_InAff_out1[0]) );
  AOI22_X1 Midori_rounds_U1047 ( .A1(reset), .A2(Midori_add_Result_Start1[53]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[53]), .ZN(
        Midori_rounds_n1899) );
  XOR2_X1 Midori_rounds_U1046 ( .A(Midori_rounds_SR_Inv_Result1[41]), .B(
        Midori_rounds_n1898), .Z(Midori_rounds_n1900) );
  OAI21_X1 Midori_rounds_U1045 ( .B1(Midori_rounds_n1897), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1896), .ZN(Midori_rounds_n845)
         );
  AOI22_X1 Midori_rounds_U1044 ( .A1(reset), .A2(Midori_add_Result_Start1[54]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result1[54]), .ZN(
        Midori_rounds_n1896) );
  XOR2_X1 Midori_rounds_U1043 ( .A(Midori_rounds_SR_Inv_Result1[42]), .B(
        Midori_rounds_n1895), .Z(Midori_rounds_n1897) );
  OAI21_X1 Midori_rounds_U1042 ( .B1(Midori_rounds_n1894), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1893), .ZN(
        Midori_rounds_sub_Sub_6_S2_InAff_out1[2]) );
  AOI22_X1 Midori_rounds_U1041 ( .A1(reset), .A2(Midori_add_Result_Start1[55]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result1[55]), .ZN(
        Midori_rounds_n1893) );
  XOR2_X1 Midori_rounds_U1040 ( .A(Midori_rounds_SR_Inv_Result1[43]), .B(
        Midori_rounds_n1892), .Z(Midori_rounds_n1894) );
  OAI21_X1 Midori_rounds_U1039 ( .B1(Midori_rounds_n1891), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1890), .ZN(
        Midori_rounds_sub_Sub_7_S1_InAff_out1[0]) );
  AOI22_X1 Midori_rounds_U1038 ( .A1(reset), .A2(Midori_add_Result_Start1[57]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result1[57]), .ZN(
        Midori_rounds_n1890) );
  XOR2_X1 Midori_rounds_U1037 ( .A(Midori_rounds_SR_Inv_Result1[21]), .B(
        Midori_rounds_n1889), .Z(Midori_rounds_n1891) );
  OAI21_X1 Midori_rounds_U1036 ( .B1(Midori_rounds_n1888), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1887), .ZN(Midori_rounds_n848)
         );
  AOI22_X1 Midori_rounds_U1035 ( .A1(reset), .A2(Midori_add_Result_Start1[58]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result1[58]), .ZN(
        Midori_rounds_n1887) );
  XOR2_X1 Midori_rounds_U1034 ( .A(Midori_rounds_SR_Inv_Result1[22]), .B(
        Midori_rounds_n1886), .Z(Midori_rounds_n1888) );
  OAI21_X1 Midori_rounds_U1033 ( .B1(Midori_rounds_n1885), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1884), .ZN(
        Midori_rounds_sub_Sub_7_S1_InAff_out1[2]) );
  AOI22_X1 Midori_rounds_U1032 ( .A1(reset), .A2(Midori_add_Result_Start1[59]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result1[59]), .ZN(
        Midori_rounds_n1884) );
  XOR2_X1 Midori_rounds_U1031 ( .A(Midori_rounds_SR_Inv_Result1[23]), .B(
        Midori_rounds_n1883), .Z(Midori_rounds_n1885) );
  OAI21_X1 Midori_rounds_U1030 ( .B1(Midori_rounds_n1882), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1881), .ZN(
        Midori_rounds_sub_Sub_7_S2_InAff_out1[0]) );
  AOI22_X1 Midori_rounds_U1029 ( .A1(reset), .A2(Midori_add_Result_Start1[61]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result1[61]), .ZN(
        Midori_rounds_n1881) );
  XOR2_X1 Midori_rounds_U1028 ( .A(Midori_rounds_SR_Inv_Result1[61]), .B(
        Midori_rounds_n1880), .Z(Midori_rounds_n1882) );
  OAI21_X1 Midori_rounds_U1027 ( .B1(Midori_rounds_n1879), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1878), .ZN(Midori_rounds_n851)
         );
  AOI22_X1 Midori_rounds_U1026 ( .A1(reset), .A2(Midori_add_Result_Start1[62]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result1[62]), .ZN(
        Midori_rounds_n1878) );
  XOR2_X1 Midori_rounds_U1025 ( .A(Midori_rounds_SR_Inv_Result1[62]), .B(
        Midori_rounds_n1877), .Z(Midori_rounds_n1879) );
  OAI21_X1 Midori_rounds_U1024 ( .B1(Midori_rounds_n1876), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1875), .ZN(
        Midori_rounds_sub_Sub_7_S2_InAff_out1[2]) );
  AOI22_X1 Midori_rounds_U1023 ( .A1(reset), .A2(Midori_add_Result_Start1[63]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result1[63]), .ZN(
        Midori_rounds_n1875) );
  XOR2_X1 Midori_rounds_U1022 ( .A(Midori_rounds_SR_Inv_Result1[63]), .B(
        Midori_rounds_n1874), .Z(Midori_rounds_n1876) );
  OAI21_X1 Midori_rounds_U1021 ( .B1(Midori_rounds_n1873), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1872), .ZN(
        Midori_rounds_sub_Sub_0_S1_InAff_out2[1]) );
  AOI22_X1 Midori_rounds_U1020 ( .A1(reset), .A2(Midori_add_Result_Start2[0]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result2[0]), .ZN(
        Midori_rounds_n1872) );
  XOR2_X1 Midori_rounds_U1019 ( .A(Midori_rounds_SR_Inv_Result2[28]), .B(
        Midori_rounds_n1871), .Z(Midori_rounds_n1873) );
  OAI21_X1 Midori_rounds_U1018 ( .B1(Midori_rounds_n1870), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1869), .ZN(
        Midori_rounds_sub_Sub_0_S1_InAff_out2[0]) );
  AOI22_X1 Midori_rounds_U1017 ( .A1(reset), .A2(Midori_add_Result_Start2[1]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result2[1]), .ZN(
        Midori_rounds_n1869) );
  XOR2_X1 Midori_rounds_U1016 ( .A(Midori_rounds_SR_Inv_Result2[29]), .B(
        Midori_rounds_n1868), .Z(Midori_rounds_n1870) );
  OAI21_X1 Midori_rounds_U1015 ( .B1(Midori_rounds_n1867), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1866), .ZN(Midori_rounds_n855)
         );
  AOI22_X1 Midori_rounds_U1014 ( .A1(reset), .A2(Midori_add_Result_Start2[2]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result2[2]), .ZN(
        Midori_rounds_n1866) );
  XOR2_X1 Midori_rounds_U1013 ( .A(Midori_rounds_SR_Inv_Result2[30]), .B(
        Midori_rounds_n1865), .Z(Midori_rounds_n1867) );
  OAI21_X1 Midori_rounds_U1012 ( .B1(Midori_rounds_n1864), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1863), .ZN(
        Midori_rounds_sub_Sub_0_S1_InAff_out2[2]) );
  AOI22_X1 Midori_rounds_U1011 ( .A1(reset), .A2(Midori_add_Result_Start2[3]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result2[3]), .ZN(
        Midori_rounds_n1863) );
  XOR2_X1 Midori_rounds_U1010 ( .A(Midori_rounds_SR_Inv_Result2[31]), .B(
        Midori_rounds_n1862), .Z(Midori_rounds_n1864) );
  OAI21_X1 Midori_rounds_U1009 ( .B1(Midori_rounds_n1861), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1860), .ZN(
        Midori_rounds_sub_Sub_0_S2_InAff_out2[1]) );
  AOI22_X1 Midori_rounds_U1008 ( .A1(reset), .A2(Midori_add_Result_Start2[4]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result2[4]), .ZN(
        Midori_rounds_n1860) );
  XOR2_X1 Midori_rounds_U1007 ( .A(Midori_rounds_SR_Inv_Result2[52]), .B(
        Midori_rounds_n1859), .Z(Midori_rounds_n1861) );
  OAI21_X1 Midori_rounds_U1006 ( .B1(Midori_rounds_n1858), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1857), .ZN(
        Midori_rounds_sub_Sub_0_S2_InAff_out2[0]) );
  AOI22_X1 Midori_rounds_U1005 ( .A1(reset), .A2(Midori_add_Result_Start2[5]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[5]), .ZN(
        Midori_rounds_n1857) );
  XOR2_X1 Midori_rounds_U1004 ( .A(Midori_rounds_SR_Inv_Result2[53]), .B(
        Midori_rounds_n1856), .Z(Midori_rounds_n1858) );
  OAI21_X1 Midori_rounds_U1003 ( .B1(Midori_rounds_n1855), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1854), .ZN(Midori_rounds_n859)
         );
  AOI22_X1 Midori_rounds_U1002 ( .A1(reset), .A2(Midori_add_Result_Start2[6]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[6]), .ZN(
        Midori_rounds_n1854) );
  XOR2_X1 Midori_rounds_U1001 ( .A(Midori_rounds_SR_Inv_Result2[54]), .B(
        Midori_rounds_n1853), .Z(Midori_rounds_n1855) );
  OAI21_X1 Midori_rounds_U1000 ( .B1(Midori_rounds_n1852), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1851), .ZN(
        Midori_rounds_sub_Sub_0_S2_InAff_out2[2]) );
  AOI22_X1 Midori_rounds_U999 ( .A1(reset), .A2(Midori_add_Result_Start2[7]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[7]), .ZN(
        Midori_rounds_n1851) );
  XOR2_X1 Midori_rounds_U998 ( .A(Midori_rounds_SR_Inv_Result2[55]), .B(
        Midori_rounds_n1850), .Z(Midori_rounds_n1852) );
  OAI21_X1 Midori_rounds_U997 ( .B1(Midori_rounds_n1849), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1848), .ZN(
        Midori_rounds_sub_Sub_1_S1_InAff_out2[1]) );
  AOI22_X1 Midori_rounds_U996 ( .A1(reset), .A2(Midori_add_Result_Start2[8]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result2[8]), .ZN(
        Midori_rounds_n1848) );
  XOR2_X1 Midori_rounds_U995 ( .A(Midori_rounds_SR_Inv_Result2[8]), .B(
        Midori_rounds_n1847), .Z(Midori_rounds_n1849) );
  OAI21_X1 Midori_rounds_U994 ( .B1(Midori_rounds_n1846), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1845), .ZN(
        Midori_rounds_sub_Sub_1_S1_InAff_out2[0]) );
  AOI22_X1 Midori_rounds_U993 ( .A1(reset), .A2(Midori_add_Result_Start2[9]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result2[9]), .ZN(
        Midori_rounds_n1845) );
  XOR2_X1 Midori_rounds_U992 ( .A(Midori_rounds_SR_Inv_Result2[9]), .B(
        Midori_rounds_n1844), .Z(Midori_rounds_n1846) );
  OAI21_X1 Midori_rounds_U991 ( .B1(Midori_rounds_n1843), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1842), .ZN(Midori_rounds_n863)
         );
  AOI22_X1 Midori_rounds_U990 ( .A1(reset), .A2(Midori_add_Result_Start2[10]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[10]), .ZN(
        Midori_rounds_n1842) );
  XOR2_X1 Midori_rounds_U989 ( .A(Midori_rounds_SR_Inv_Result2[10]), .B(
        Midori_rounds_n1841), .Z(Midori_rounds_n1843) );
  OAI21_X1 Midori_rounds_U988 ( .B1(Midori_rounds_n1840), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1839), .ZN(
        Midori_rounds_sub_Sub_1_S1_InAff_out2[2]) );
  AOI22_X1 Midori_rounds_U987 ( .A1(reset), .A2(Midori_add_Result_Start2[11]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[11]), .ZN(
        Midori_rounds_n1839) );
  XOR2_X1 Midori_rounds_U986 ( .A(Midori_rounds_SR_Inv_Result2[11]), .B(
        Midori_rounds_n1838), .Z(Midori_rounds_n1840) );
  OAI21_X1 Midori_rounds_U985 ( .B1(Midori_rounds_n1837), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1836), .ZN(
        Midori_rounds_sub_Sub_1_S2_InAff_out2[1]) );
  AOI22_X1 Midori_rounds_U984 ( .A1(reset), .A2(Midori_add_Result_Start2[12]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[12]), .ZN(
        Midori_rounds_n1836) );
  XOR2_X1 Midori_rounds_U983 ( .A(Midori_rounds_SR_Inv_Result2[32]), .B(
        Midori_rounds_n1835), .Z(Midori_rounds_n1837) );
  OAI21_X1 Midori_rounds_U982 ( .B1(Midori_rounds_n1834), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1833), .ZN(
        Midori_rounds_sub_Sub_1_S2_InAff_out2[0]) );
  AOI22_X1 Midori_rounds_U981 ( .A1(reset), .A2(Midori_add_Result_Start2[13]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result2[13]), .ZN(
        Midori_rounds_n1833) );
  XOR2_X1 Midori_rounds_U980 ( .A(Midori_rounds_SR_Inv_Result2[33]), .B(
        Midori_rounds_n1832), .Z(Midori_rounds_n1834) );
  OAI21_X1 Midori_rounds_U979 ( .B1(Midori_rounds_n1831), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1830), .ZN(Midori_rounds_n867)
         );
  AOI22_X1 Midori_rounds_U978 ( .A1(reset), .A2(Midori_add_Result_Start2[14]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result2[14]), .ZN(
        Midori_rounds_n1830) );
  XOR2_X1 Midori_rounds_U977 ( .A(Midori_rounds_SR_Inv_Result2[34]), .B(
        Midori_rounds_n1829), .Z(Midori_rounds_n1831) );
  OAI21_X1 Midori_rounds_U976 ( .B1(Midori_rounds_n1828), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1827), .ZN(
        Midori_rounds_sub_Sub_1_S2_InAff_out2[2]) );
  AOI22_X1 Midori_rounds_U975 ( .A1(reset), .A2(Midori_add_Result_Start2[15]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result2[15]), .ZN(
        Midori_rounds_n1827) );
  XOR2_X1 Midori_rounds_U974 ( .A(Midori_rounds_SR_Inv_Result2[35]), .B(
        Midori_rounds_n1826), .Z(Midori_rounds_n1828) );
  OAI21_X1 Midori_rounds_U973 ( .B1(Midori_rounds_n1825), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1824), .ZN(
        Midori_rounds_sub_Sub_2_S1_InAff_out2[1]) );
  AOI22_X1 Midori_rounds_U972 ( .A1(reset), .A2(Midori_add_Result_Start2[16]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result2[16]), .ZN(
        Midori_rounds_n1824) );
  XOR2_X1 Midori_rounds_U971 ( .A(Midori_rounds_SR_Inv_Result2[36]), .B(
        Midori_rounds_n1823), .Z(Midori_rounds_n1825) );
  OAI21_X1 Midori_rounds_U970 ( .B1(Midori_rounds_n1822), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1821), .ZN(
        Midori_rounds_sub_Sub_2_S1_InAff_out2[0]) );
  AOI22_X1 Midori_rounds_U969 ( .A1(reset), .A2(Midori_add_Result_Start2[17]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result2[17]), .ZN(
        Midori_rounds_n1821) );
  XOR2_X1 Midori_rounds_U968 ( .A(Midori_rounds_SR_Inv_Result2[37]), .B(
        Midori_rounds_n1820), .Z(Midori_rounds_n1822) );
  OAI21_X1 Midori_rounds_U967 ( .B1(Midori_rounds_n1819), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1818), .ZN(Midori_rounds_n871)
         );
  AOI22_X1 Midori_rounds_U966 ( .A1(reset), .A2(Midori_add_Result_Start2[18]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result2[18]), .ZN(
        Midori_rounds_n1818) );
  XOR2_X1 Midori_rounds_U965 ( .A(Midori_rounds_SR_Inv_Result2[38]), .B(
        Midori_rounds_n1817), .Z(Midori_rounds_n1819) );
  OAI21_X1 Midori_rounds_U964 ( .B1(Midori_rounds_n1816), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1815), .ZN(
        Midori_rounds_sub_Sub_2_S1_InAff_out2[2]) );
  AOI22_X1 Midori_rounds_U963 ( .A1(reset), .A2(Midori_add_Result_Start2[19]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result2[19]), .ZN(
        Midori_rounds_n1815) );
  XOR2_X1 Midori_rounds_U962 ( .A(Midori_rounds_SR_Inv_Result2[39]), .B(
        Midori_rounds_n1814), .Z(Midori_rounds_n1816) );
  OAI21_X1 Midori_rounds_U961 ( .B1(Midori_rounds_n1813), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1812), .ZN(
        Midori_rounds_sub_Sub_2_S2_InAff_out2[1]) );
  AOI22_X1 Midori_rounds_U960 ( .A1(reset), .A2(Midori_add_Result_Start2[20]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result2[20]), .ZN(
        Midori_rounds_n1812) );
  XOR2_X1 Midori_rounds_U959 ( .A(Midori_rounds_SR_Inv_Result2[12]), .B(
        Midori_rounds_n1811), .Z(Midori_rounds_n1813) );
  OAI21_X1 Midori_rounds_U958 ( .B1(Midori_rounds_n1810), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1809), .ZN(
        Midori_rounds_sub_Sub_2_S2_InAff_out2[0]) );
  AOI22_X1 Midori_rounds_U957 ( .A1(reset), .A2(Midori_add_Result_Start2[21]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result2[21]), .ZN(
        Midori_rounds_n1809) );
  XOR2_X1 Midori_rounds_U956 ( .A(Midori_rounds_SR_Inv_Result2[13]), .B(
        Midori_rounds_n1808), .Z(Midori_rounds_n1810) );
  OAI21_X1 Midori_rounds_U955 ( .B1(Midori_rounds_n1807), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1806), .ZN(Midori_rounds_n875)
         );
  AOI22_X1 Midori_rounds_U954 ( .A1(reset), .A2(Midori_add_Result_Start2[22]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result2[22]), .ZN(
        Midori_rounds_n1806) );
  XOR2_X1 Midori_rounds_U953 ( .A(Midori_rounds_SR_Inv_Result2[14]), .B(
        Midori_rounds_n1805), .Z(Midori_rounds_n1807) );
  OAI21_X1 Midori_rounds_U952 ( .B1(Midori_rounds_n1804), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1803), .ZN(
        Midori_rounds_sub_Sub_2_S2_InAff_out2[2]) );
  AOI22_X1 Midori_rounds_U951 ( .A1(reset), .A2(Midori_add_Result_Start2[23]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[23]), .ZN(
        Midori_rounds_n1803) );
  XOR2_X1 Midori_rounds_U950 ( .A(Midori_rounds_SR_Inv_Result2[15]), .B(
        Midori_rounds_n1802), .Z(Midori_rounds_n1804) );
  OAI21_X1 Midori_rounds_U949 ( .B1(Midori_rounds_n1801), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1800), .ZN(
        Midori_rounds_sub_Sub_3_S1_InAff_out2[1]) );
  AOI22_X1 Midori_rounds_U948 ( .A1(reset), .A2(Midori_add_Result_Start2[24]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[24]), .ZN(
        Midori_rounds_n1800) );
  XOR2_X1 Midori_rounds_U947 ( .A(Midori_rounds_SR_Inv_Result2[48]), .B(
        Midori_rounds_n1799), .Z(Midori_rounds_n1801) );
  OAI21_X1 Midori_rounds_U946 ( .B1(Midori_rounds_n1798), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1797), .ZN(
        Midori_rounds_sub_Sub_3_S1_InAff_out2[0]) );
  AOI22_X1 Midori_rounds_U945 ( .A1(reset), .A2(Midori_add_Result_Start2[25]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[25]), .ZN(
        Midori_rounds_n1797) );
  XOR2_X1 Midori_rounds_U944 ( .A(Midori_rounds_SR_Inv_Result2[49]), .B(
        Midori_rounds_n1796), .Z(Midori_rounds_n1798) );
  OAI21_X1 Midori_rounds_U943 ( .B1(Midori_rounds_n1795), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1794), .ZN(Midori_rounds_n879)
         );
  AOI22_X1 Midori_rounds_U942 ( .A1(reset), .A2(Midori_add_Result_Start2[26]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result2[26]), .ZN(
        Midori_rounds_n1794) );
  XOR2_X1 Midori_rounds_U941 ( .A(Midori_rounds_SR_Inv_Result2[50]), .B(
        Midori_rounds_n1793), .Z(Midori_rounds_n1795) );
  OAI21_X1 Midori_rounds_U940 ( .B1(Midori_rounds_n1792), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1791), .ZN(
        Midori_rounds_sub_Sub_3_S1_InAff_out2[2]) );
  AOI22_X1 Midori_rounds_U939 ( .A1(reset), .A2(Midori_add_Result_Start2[27]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result2[27]), .ZN(
        Midori_rounds_n1791) );
  XOR2_X1 Midori_rounds_U938 ( .A(Midori_rounds_SR_Inv_Result2[51]), .B(
        Midori_rounds_n1790), .Z(Midori_rounds_n1792) );
  OAI21_X1 Midori_rounds_U937 ( .B1(Midori_rounds_n1789), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1788), .ZN(
        Midori_rounds_sub_Sub_3_S2_InAff_out2[1]) );
  AOI22_X1 Midori_rounds_U936 ( .A1(reset), .A2(Midori_add_Result_Start2[28]), 
        .B1(Midori_rounds_n1259), .B2(Midori_rounds_SR_Inv_Result2[28]), .ZN(
        Midori_rounds_n1788) );
  XOR2_X1 Midori_rounds_U935 ( .A(Midori_rounds_SR_Inv_Result2[24]), .B(
        Midori_rounds_n1787), .Z(Midori_rounds_n1789) );
  OAI21_X1 Midori_rounds_U934 ( .B1(Midori_rounds_n1786), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1785), .ZN(
        Midori_rounds_sub_Sub_3_S2_InAff_out2[0]) );
  AOI22_X1 Midori_rounds_U933 ( .A1(reset), .A2(Midori_add_Result_Start2[29]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result2[29]), .ZN(
        Midori_rounds_n1785) );
  XOR2_X1 Midori_rounds_U932 ( .A(Midori_rounds_SR_Inv_Result2[25]), .B(
        Midori_rounds_n1784), .Z(Midori_rounds_n1786) );
  OAI21_X1 Midori_rounds_U931 ( .B1(Midori_rounds_n1783), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1782), .ZN(Midori_rounds_n883)
         );
  AOI22_X1 Midori_rounds_U930 ( .A1(reset), .A2(Midori_add_Result_Start2[30]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result2[30]), .ZN(
        Midori_rounds_n1782) );
  XOR2_X1 Midori_rounds_U929 ( .A(Midori_rounds_SR_Inv_Result2[26]), .B(
        Midori_rounds_n1781), .Z(Midori_rounds_n1783) );
  OAI21_X1 Midori_rounds_U928 ( .B1(Midori_rounds_n1780), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1779), .ZN(
        Midori_rounds_sub_Sub_3_S2_InAff_out2[2]) );
  AOI22_X1 Midori_rounds_U927 ( .A1(reset), .A2(Midori_add_Result_Start2[31]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[31]), .ZN(
        Midori_rounds_n1779) );
  XOR2_X1 Midori_rounds_U926 ( .A(Midori_rounds_SR_Inv_Result2[27]), .B(
        Midori_rounds_n1778), .Z(Midori_rounds_n1780) );
  OAI21_X1 Midori_rounds_U925 ( .B1(Midori_rounds_n1777), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1776), .ZN(
        Midori_rounds_sub_Sub_4_S1_InAff_out2[1]) );
  AOI22_X1 Midori_rounds_U924 ( .A1(reset), .A2(Midori_add_Result_Start2[32]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[32]), .ZN(
        Midori_rounds_n1776) );
  XOR2_X1 Midori_rounds_U923 ( .A(Midori_rounds_SR_Inv_Result2[56]), .B(
        Midori_rounds_n1775), .Z(Midori_rounds_n1777) );
  OAI21_X1 Midori_rounds_U922 ( .B1(Midori_rounds_n1774), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1773), .ZN(
        Midori_rounds_sub_Sub_4_S1_InAff_out2[0]) );
  AOI22_X1 Midori_rounds_U921 ( .A1(reset), .A2(Midori_add_Result_Start2[33]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[33]), .ZN(
        Midori_rounds_n1773) );
  XOR2_X1 Midori_rounds_U920 ( .A(Midori_rounds_SR_Inv_Result2[57]), .B(
        Midori_rounds_n1772), .Z(Midori_rounds_n1774) );
  OAI21_X1 Midori_rounds_U919 ( .B1(Midori_rounds_n1771), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1770), .ZN(Midori_rounds_n887)
         );
  AOI22_X1 Midori_rounds_U918 ( .A1(reset), .A2(Midori_add_Result_Start2[34]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[34]), .ZN(
        Midori_rounds_n1770) );
  XOR2_X1 Midori_rounds_U917 ( .A(Midori_rounds_SR_Inv_Result2[58]), .B(
        Midori_rounds_n1769), .Z(Midori_rounds_n1771) );
  OAI21_X1 Midori_rounds_U916 ( .B1(Midori_rounds_n1768), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1767), .ZN(
        Midori_rounds_sub_Sub_4_S1_InAff_out2[2]) );
  AOI22_X1 Midori_rounds_U915 ( .A1(reset), .A2(Midori_add_Result_Start2[35]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[35]), .ZN(
        Midori_rounds_n1767) );
  XOR2_X1 Midori_rounds_U914 ( .A(Midori_rounds_SR_Inv_Result2[59]), .B(
        Midori_rounds_n1766), .Z(Midori_rounds_n1768) );
  OAI21_X1 Midori_rounds_U913 ( .B1(Midori_rounds_n1765), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1764), .ZN(
        Midori_rounds_sub_Sub_4_S2_InAff_out2[1]) );
  AOI22_X1 Midori_rounds_U912 ( .A1(reset), .A2(Midori_add_Result_Start2[36]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[36]), .ZN(
        Midori_rounds_n1764) );
  XOR2_X1 Midori_rounds_U911 ( .A(Midori_rounds_SR_Inv_Result2[16]), .B(
        Midori_rounds_n1763), .Z(Midori_rounds_n1765) );
  OAI21_X1 Midori_rounds_U910 ( .B1(Midori_rounds_n1762), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1761), .ZN(
        Midori_rounds_sub_Sub_4_S2_InAff_out2[0]) );
  AOI22_X1 Midori_rounds_U909 ( .A1(reset), .A2(Midori_add_Result_Start2[37]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[37]), .ZN(
        Midori_rounds_n1761) );
  XOR2_X1 Midori_rounds_U908 ( .A(Midori_rounds_SR_Inv_Result2[17]), .B(
        Midori_rounds_n1760), .Z(Midori_rounds_n1762) );
  OAI21_X1 Midori_rounds_U907 ( .B1(Midori_rounds_n1759), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1758), .ZN(Midori_rounds_n891)
         );
  AOI22_X1 Midori_rounds_U906 ( .A1(reset), .A2(Midori_add_Result_Start2[38]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[38]), .ZN(
        Midori_rounds_n1758) );
  XOR2_X1 Midori_rounds_U905 ( .A(Midori_rounds_SR_Inv_Result2[18]), .B(
        Midori_rounds_n1757), .Z(Midori_rounds_n1759) );
  OAI21_X1 Midori_rounds_U904 ( .B1(Midori_rounds_n1756), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1755), .ZN(
        Midori_rounds_sub_Sub_4_S2_InAff_out2[2]) );
  AOI22_X1 Midori_rounds_U903 ( .A1(reset), .A2(Midori_add_Result_Start2[39]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[39]), .ZN(
        Midori_rounds_n1755) );
  XOR2_X1 Midori_rounds_U902 ( .A(Midori_rounds_SR_Inv_Result2[19]), .B(
        Midori_rounds_n1754), .Z(Midori_rounds_n1756) );
  OAI21_X1 Midori_rounds_U901 ( .B1(Midori_rounds_n1753), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1752), .ZN(
        Midori_rounds_sub_Sub_5_S1_InAff_out2[1]) );
  AOI22_X1 Midori_rounds_U900 ( .A1(reset), .A2(Midori_add_Result_Start2[40]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[40]), .ZN(
        Midori_rounds_n1752) );
  XOR2_X1 Midori_rounds_U899 ( .A(Midori_rounds_SR_Inv_Result2[44]), .B(
        Midori_rounds_n1751), .Z(Midori_rounds_n1753) );
  OAI21_X1 Midori_rounds_U898 ( .B1(Midori_rounds_n1750), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1749), .ZN(
        Midori_rounds_sub_Sub_5_S1_InAff_out2[0]) );
  AOI22_X1 Midori_rounds_U897 ( .A1(reset), .A2(Midori_add_Result_Start2[41]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[41]), .ZN(
        Midori_rounds_n1749) );
  XOR2_X1 Midori_rounds_U896 ( .A(Midori_rounds_SR_Inv_Result2[45]), .B(
        Midori_rounds_n1748), .Z(Midori_rounds_n1750) );
  OAI21_X1 Midori_rounds_U895 ( .B1(Midori_rounds_n1747), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1746), .ZN(Midori_rounds_n895)
         );
  AOI22_X1 Midori_rounds_U894 ( .A1(reset), .A2(Midori_add_Result_Start2[42]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[42]), .ZN(
        Midori_rounds_n1746) );
  XOR2_X1 Midori_rounds_U893 ( .A(Midori_rounds_SR_Inv_Result2[46]), .B(
        Midori_rounds_n1745), .Z(Midori_rounds_n1747) );
  OAI21_X1 Midori_rounds_U892 ( .B1(Midori_rounds_n1744), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1743), .ZN(
        Midori_rounds_sub_Sub_5_S1_InAff_out2[2]) );
  AOI22_X1 Midori_rounds_U891 ( .A1(reset), .A2(Midori_add_Result_Start2[43]), 
        .B1(Midori_rounds_n1258), .B2(Midori_rounds_SR_Inv_Result2[43]), .ZN(
        Midori_rounds_n1743) );
  XOR2_X1 Midori_rounds_U890 ( .A(Midori_rounds_SR_Inv_Result2[47]), .B(
        Midori_rounds_n1742), .Z(Midori_rounds_n1744) );
  OAI21_X1 Midori_rounds_U889 ( .B1(Midori_rounds_n1741), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1740), .ZN(
        Midori_rounds_sub_Sub_5_S2_InAff_out2[1]) );
  AOI22_X1 Midori_rounds_U888 ( .A1(reset), .A2(Midori_add_Result_Start2[44]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[44]), .ZN(
        Midori_rounds_n1740) );
  XOR2_X1 Midori_rounds_U887 ( .A(Midori_rounds_SR_Inv_Result2[4]), .B(
        Midori_rounds_n1739), .Z(Midori_rounds_n1741) );
  OAI21_X1 Midori_rounds_U886 ( .B1(Midori_rounds_n1738), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1737), .ZN(
        Midori_rounds_sub_Sub_5_S2_InAff_out2[0]) );
  AOI22_X1 Midori_rounds_U885 ( .A1(reset), .A2(Midori_add_Result_Start2[45]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[45]), .ZN(
        Midori_rounds_n1737) );
  XOR2_X1 Midori_rounds_U884 ( .A(Midori_rounds_SR_Inv_Result2[5]), .B(
        Midori_rounds_n1736), .Z(Midori_rounds_n1738) );
  OAI21_X1 Midori_rounds_U883 ( .B1(Midori_rounds_n1735), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1734), .ZN(Midori_rounds_n899)
         );
  AOI22_X1 Midori_rounds_U882 ( .A1(reset), .A2(Midori_add_Result_Start2[46]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[46]), .ZN(
        Midori_rounds_n1734) );
  XOR2_X1 Midori_rounds_U881 ( .A(Midori_rounds_SR_Inv_Result2[6]), .B(
        Midori_rounds_n1733), .Z(Midori_rounds_n1735) );
  OAI21_X1 Midori_rounds_U880 ( .B1(Midori_rounds_n1732), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1731), .ZN(
        Midori_rounds_sub_Sub_5_S2_InAff_out2[2]) );
  AOI22_X1 Midori_rounds_U879 ( .A1(reset), .A2(Midori_add_Result_Start2[47]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[47]), .ZN(
        Midori_rounds_n1731) );
  XOR2_X1 Midori_rounds_U878 ( .A(Midori_rounds_SR_Inv_Result2[7]), .B(
        Midori_rounds_n1730), .Z(Midori_rounds_n1732) );
  OAI21_X1 Midori_rounds_U877 ( .B1(Midori_rounds_n1729), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1728), .ZN(
        Midori_rounds_sub_Sub_6_S1_InAff_out2[1]) );
  AOI22_X1 Midori_rounds_U876 ( .A1(reset), .A2(Midori_add_Result_Start2[48]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[48]), .ZN(
        Midori_rounds_n1728) );
  XOR2_X1 Midori_rounds_U875 ( .A(Midori_rounds_SR_Inv_Result2[0]), .B(
        Midori_rounds_n1727), .Z(Midori_rounds_n1729) );
  OAI21_X1 Midori_rounds_U874 ( .B1(Midori_rounds_n1726), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1725), .ZN(
        Midori_rounds_sub_Sub_6_S1_InAff_out2[0]) );
  AOI22_X1 Midori_rounds_U873 ( .A1(reset), .A2(Midori_add_Result_Start2[49]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[49]), .ZN(
        Midori_rounds_n1725) );
  XOR2_X1 Midori_rounds_U872 ( .A(Midori_rounds_SR_Inv_Result2[1]), .B(
        Midori_rounds_n1724), .Z(Midori_rounds_n1726) );
  OAI21_X1 Midori_rounds_U871 ( .B1(Midori_rounds_n1723), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1722), .ZN(Midori_rounds_n903)
         );
  AOI22_X1 Midori_rounds_U870 ( .A1(reset), .A2(Midori_add_Result_Start2[50]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[50]), .ZN(
        Midori_rounds_n1722) );
  XOR2_X1 Midori_rounds_U869 ( .A(Midori_rounds_SR_Inv_Result2[2]), .B(
        Midori_rounds_n1721), .Z(Midori_rounds_n1723) );
  OAI21_X1 Midori_rounds_U868 ( .B1(Midori_rounds_n1720), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1719), .ZN(
        Midori_rounds_sub_Sub_6_S1_InAff_out2[2]) );
  AOI22_X1 Midori_rounds_U867 ( .A1(reset), .A2(Midori_add_Result_Start2[51]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[51]), .ZN(
        Midori_rounds_n1719) );
  XOR2_X1 Midori_rounds_U866 ( .A(Midori_rounds_SR_Inv_Result2[3]), .B(
        Midori_rounds_n1718), .Z(Midori_rounds_n1720) );
  OAI21_X1 Midori_rounds_U865 ( .B1(Midori_rounds_n1717), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1716), .ZN(
        Midori_rounds_sub_Sub_6_S2_InAff_out2[1]) );
  AOI22_X1 Midori_rounds_U864 ( .A1(reset), .A2(Midori_add_Result_Start2[52]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[52]), .ZN(
        Midori_rounds_n1716) );
  XOR2_X1 Midori_rounds_U863 ( .A(Midori_rounds_SR_Inv_Result2[40]), .B(
        Midori_rounds_n1715), .Z(Midori_rounds_n1717) );
  OAI21_X1 Midori_rounds_U862 ( .B1(Midori_rounds_n1714), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1713), .ZN(
        Midori_rounds_sub_Sub_6_S2_InAff_out2[0]) );
  AOI22_X1 Midori_rounds_U861 ( .A1(reset), .A2(Midori_add_Result_Start2[53]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[53]), .ZN(
        Midori_rounds_n1713) );
  XOR2_X1 Midori_rounds_U860 ( .A(Midori_rounds_SR_Inv_Result2[41]), .B(
        Midori_rounds_n1712), .Z(Midori_rounds_n1714) );
  OAI21_X1 Midori_rounds_U859 ( .B1(Midori_rounds_n1711), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1710), .ZN(Midori_rounds_n907)
         );
  AOI22_X1 Midori_rounds_U858 ( .A1(reset), .A2(Midori_add_Result_Start2[54]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[54]), .ZN(
        Midori_rounds_n1710) );
  XOR2_X1 Midori_rounds_U857 ( .A(Midori_rounds_SR_Inv_Result2[42]), .B(
        Midori_rounds_n1709), .Z(Midori_rounds_n1711) );
  OAI21_X1 Midori_rounds_U856 ( .B1(Midori_rounds_n1708), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1707), .ZN(
        Midori_rounds_sub_Sub_6_S2_InAff_out2[2]) );
  AOI22_X1 Midori_rounds_U855 ( .A1(reset), .A2(Midori_add_Result_Start2[55]), 
        .B1(Midori_rounds_n1257), .B2(Midori_rounds_SR_Inv_Result2[55]), .ZN(
        Midori_rounds_n1707) );
  XOR2_X1 Midori_rounds_U854 ( .A(Midori_rounds_SR_Inv_Result2[43]), .B(
        Midori_rounds_n1706), .Z(Midori_rounds_n1708) );
  OAI21_X1 Midori_rounds_U853 ( .B1(Midori_rounds_n1705), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1704), .ZN(
        Midori_rounds_sub_Sub_7_S1_InAff_out2[1]) );
  AOI22_X1 Midori_rounds_U852 ( .A1(reset), .A2(Midori_add_Result_Start2[56]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[56]), .ZN(
        Midori_rounds_n1704) );
  XOR2_X1 Midori_rounds_U851 ( .A(Midori_rounds_SR_Inv_Result2[20]), .B(
        Midori_rounds_n1703), .Z(Midori_rounds_n1705) );
  OAI21_X1 Midori_rounds_U850 ( .B1(Midori_rounds_n1702), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1701), .ZN(
        Midori_rounds_sub_Sub_7_S1_InAff_out2[0]) );
  AOI22_X1 Midori_rounds_U849 ( .A1(reset), .A2(Midori_add_Result_Start2[57]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[57]), .ZN(
        Midori_rounds_n1701) );
  XOR2_X1 Midori_rounds_U848 ( .A(Midori_rounds_SR_Inv_Result2[21]), .B(
        Midori_rounds_n1700), .Z(Midori_rounds_n1702) );
  OAI21_X1 Midori_rounds_U847 ( .B1(Midori_rounds_n1699), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1698), .ZN(Midori_rounds_n911)
         );
  AOI22_X1 Midori_rounds_U846 ( .A1(reset), .A2(Midori_add_Result_Start2[58]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[58]), .ZN(
        Midori_rounds_n1698) );
  XOR2_X1 Midori_rounds_U845 ( .A(Midori_rounds_SR_Inv_Result2[22]), .B(
        Midori_rounds_n1697), .Z(Midori_rounds_n1699) );
  OAI21_X1 Midori_rounds_U844 ( .B1(Midori_rounds_n1696), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1695), .ZN(
        Midori_rounds_sub_Sub_7_S1_InAff_out2[2]) );
  AOI22_X1 Midori_rounds_U843 ( .A1(reset), .A2(Midori_add_Result_Start2[59]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[59]), .ZN(
        Midori_rounds_n1695) );
  XOR2_X1 Midori_rounds_U842 ( .A(Midori_rounds_SR_Inv_Result2[23]), .B(
        Midori_rounds_n1694), .Z(Midori_rounds_n1696) );
  OAI21_X1 Midori_rounds_U841 ( .B1(Midori_rounds_n1693), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1692), .ZN(
        Midori_rounds_sub_Sub_7_S2_InAff_out2[1]) );
  AOI22_X1 Midori_rounds_U840 ( .A1(reset), .A2(Midori_add_Result_Start2[60]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[60]), .ZN(
        Midori_rounds_n1692) );
  XOR2_X1 Midori_rounds_U839 ( .A(Midori_rounds_SR_Inv_Result2[60]), .B(
        Midori_rounds_n1691), .Z(Midori_rounds_n1693) );
  OAI21_X1 Midori_rounds_U838 ( .B1(Midori_rounds_n1690), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1689), .ZN(
        Midori_rounds_sub_Sub_7_S2_InAff_out2[0]) );
  AOI22_X1 Midori_rounds_U837 ( .A1(reset), .A2(Midori_add_Result_Start2[61]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[61]), .ZN(
        Midori_rounds_n1689) );
  XOR2_X1 Midori_rounds_U836 ( .A(Midori_rounds_SR_Inv_Result2[61]), .B(
        Midori_rounds_n1688), .Z(Midori_rounds_n1690) );
  OAI21_X1 Midori_rounds_U835 ( .B1(Midori_rounds_n1687), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1686), .ZN(Midori_rounds_n915)
         );
  AOI22_X1 Midori_rounds_U834 ( .A1(reset), .A2(Midori_add_Result_Start2[62]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[62]), .ZN(
        Midori_rounds_n1686) );
  XOR2_X1 Midori_rounds_U833 ( .A(Midori_rounds_SR_Inv_Result2[62]), .B(
        Midori_rounds_n1685), .Z(Midori_rounds_n1687) );
  OAI21_X1 Midori_rounds_U832 ( .B1(Midori_rounds_n1684), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1683), .ZN(
        Midori_rounds_sub_Sub_7_S2_InAff_out2[2]) );
  AOI22_X1 Midori_rounds_U831 ( .A1(reset), .A2(Midori_add_Result_Start2[63]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result2[63]), .ZN(
        Midori_rounds_n1683) );
  XOR2_X1 Midori_rounds_U830 ( .A(Midori_rounds_SR_Inv_Result2[63]), .B(
        Midori_rounds_n1682), .Z(Midori_rounds_n1684) );
  OAI21_X1 Midori_rounds_U829 ( .B1(Midori_rounds_n1681), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1680), .ZN(
        Midori_rounds_sub_Sub_0_S1_InAff_out3[1]) );
  AOI22_X1 Midori_rounds_U828 ( .A1(reset), .A2(Midori_add_Result_Start3[0]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result3[0]), .ZN(
        Midori_rounds_n1680) );
  XOR2_X1 Midori_rounds_U827 ( .A(Midori_rounds_SR_Inv_Result3[28]), .B(
        Midori_rounds_n1679), .Z(Midori_rounds_n1681) );
  OAI21_X1 Midori_rounds_U826 ( .B1(Midori_rounds_n1678), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1677), .ZN(
        Midori_rounds_sub_Sub_0_S1_InAff_out3[0]) );
  AOI22_X1 Midori_rounds_U825 ( .A1(reset), .A2(Midori_add_Result_Start3[1]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result3[1]), .ZN(
        Midori_rounds_n1677) );
  XOR2_X1 Midori_rounds_U824 ( .A(Midori_rounds_SR_Inv_Result3[29]), .B(
        Midori_rounds_n1676), .Z(Midori_rounds_n1678) );
  OAI21_X1 Midori_rounds_U823 ( .B1(Midori_rounds_n1675), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1674), .ZN(Midori_rounds_n919)
         );
  AOI22_X1 Midori_rounds_U822 ( .A1(reset), .A2(Midori_add_Result_Start3[2]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result3[2]), .ZN(
        Midori_rounds_n1674) );
  XOR2_X1 Midori_rounds_U821 ( .A(Midori_rounds_SR_Inv_Result3[30]), .B(
        Midori_rounds_n1673), .Z(Midori_rounds_n1675) );
  OAI21_X1 Midori_rounds_U820 ( .B1(Midori_rounds_n1672), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1671), .ZN(
        Midori_rounds_sub_Sub_0_S1_InAff_out3[2]) );
  AOI22_X1 Midori_rounds_U819 ( .A1(reset), .A2(Midori_add_Result_Start3[3]), 
        .B1(Midori_rounds_n1256), .B2(Midori_rounds_SR_Inv_Result3[3]), .ZN(
        Midori_rounds_n1671) );
  XOR2_X1 Midori_rounds_U818 ( .A(Midori_rounds_SR_Inv_Result3[31]), .B(
        Midori_rounds_n1670), .Z(Midori_rounds_n1672) );
  OAI21_X1 Midori_rounds_U817 ( .B1(Midori_rounds_n1669), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1668), .ZN(
        Midori_rounds_sub_Sub_0_S2_InAff_out3[1]) );
  AOI22_X1 Midori_rounds_U816 ( .A1(reset), .A2(Midori_add_Result_Start3[4]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[4]), .ZN(
        Midori_rounds_n1668) );
  XOR2_X1 Midori_rounds_U815 ( .A(Midori_rounds_SR_Inv_Result3[52]), .B(
        Midori_rounds_n1667), .Z(Midori_rounds_n1669) );
  OAI21_X1 Midori_rounds_U814 ( .B1(Midori_rounds_n1666), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1665), .ZN(
        Midori_rounds_sub_Sub_0_S2_InAff_out3[0]) );
  AOI22_X1 Midori_rounds_U813 ( .A1(reset), .A2(Midori_add_Result_Start3[5]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[5]), .ZN(
        Midori_rounds_n1665) );
  XOR2_X1 Midori_rounds_U812 ( .A(Midori_rounds_SR_Inv_Result3[53]), .B(
        Midori_rounds_n1664), .Z(Midori_rounds_n1666) );
  OAI21_X1 Midori_rounds_U811 ( .B1(Midori_rounds_n1663), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1662), .ZN(Midori_rounds_n923)
         );
  AOI22_X1 Midori_rounds_U810 ( .A1(reset), .A2(Midori_add_Result_Start3[6]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[6]), .ZN(
        Midori_rounds_n1662) );
  XOR2_X1 Midori_rounds_U809 ( .A(Midori_rounds_SR_Inv_Result3[54]), .B(
        Midori_rounds_n1661), .Z(Midori_rounds_n1663) );
  OAI21_X1 Midori_rounds_U808 ( .B1(Midori_rounds_n1660), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1659), .ZN(
        Midori_rounds_sub_Sub_0_S2_InAff_out3[2]) );
  AOI22_X1 Midori_rounds_U807 ( .A1(reset), .A2(Midori_add_Result_Start3[7]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[7]), .ZN(
        Midori_rounds_n1659) );
  XOR2_X1 Midori_rounds_U806 ( .A(Midori_rounds_SR_Inv_Result3[55]), .B(
        Midori_rounds_n1658), .Z(Midori_rounds_n1660) );
  OAI21_X1 Midori_rounds_U805 ( .B1(Midori_rounds_n1657), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1656), .ZN(
        Midori_rounds_sub_Sub_1_S1_InAff_out3[1]) );
  AOI22_X1 Midori_rounds_U804 ( .A1(reset), .A2(Midori_add_Result_Start3[8]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[8]), .ZN(
        Midori_rounds_n1656) );
  XOR2_X1 Midori_rounds_U803 ( .A(Midori_rounds_SR_Inv_Result3[8]), .B(
        Midori_rounds_n1655), .Z(Midori_rounds_n1657) );
  OAI21_X1 Midori_rounds_U802 ( .B1(Midori_rounds_n1654), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1653), .ZN(
        Midori_rounds_sub_Sub_1_S1_InAff_out3[0]) );
  AOI22_X1 Midori_rounds_U801 ( .A1(reset), .A2(Midori_add_Result_Start3[9]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[9]), .ZN(
        Midori_rounds_n1653) );
  XOR2_X1 Midori_rounds_U800 ( .A(Midori_rounds_SR_Inv_Result3[9]), .B(
        Midori_rounds_n1652), .Z(Midori_rounds_n1654) );
  OAI21_X1 Midori_rounds_U799 ( .B1(Midori_rounds_n1651), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1650), .ZN(Midori_rounds_n927)
         );
  AOI22_X1 Midori_rounds_U798 ( .A1(reset), .A2(Midori_add_Result_Start3[10]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[10]), .ZN(
        Midori_rounds_n1650) );
  XOR2_X1 Midori_rounds_U797 ( .A(Midori_rounds_SR_Inv_Result3[10]), .B(
        Midori_rounds_n1649), .Z(Midori_rounds_n1651) );
  OAI21_X1 Midori_rounds_U796 ( .B1(Midori_rounds_n1648), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1647), .ZN(
        Midori_rounds_sub_Sub_1_S1_InAff_out3[2]) );
  AOI22_X1 Midori_rounds_U795 ( .A1(reset), .A2(Midori_add_Result_Start3[11]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[11]), .ZN(
        Midori_rounds_n1647) );
  XOR2_X1 Midori_rounds_U794 ( .A(Midori_rounds_SR_Inv_Result3[11]), .B(
        Midori_rounds_n1646), .Z(Midori_rounds_n1648) );
  OAI21_X1 Midori_rounds_U793 ( .B1(Midori_rounds_n1645), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1644), .ZN(
        Midori_rounds_sub_Sub_1_S2_InAff_out3[1]) );
  AOI22_X1 Midori_rounds_U792 ( .A1(reset), .A2(Midori_add_Result_Start3[12]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[12]), .ZN(
        Midori_rounds_n1644) );
  XOR2_X1 Midori_rounds_U791 ( .A(Midori_rounds_SR_Inv_Result3[32]), .B(
        Midori_rounds_n1643), .Z(Midori_rounds_n1645) );
  OAI21_X1 Midori_rounds_U790 ( .B1(Midori_rounds_n1642), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1641), .ZN(
        Midori_rounds_sub_Sub_1_S2_InAff_out3[0]) );
  AOI22_X1 Midori_rounds_U789 ( .A1(reset), .A2(Midori_add_Result_Start3[13]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[13]), .ZN(
        Midori_rounds_n1641) );
  XOR2_X1 Midori_rounds_U788 ( .A(Midori_rounds_SR_Inv_Result3[33]), .B(
        Midori_rounds_n1640), .Z(Midori_rounds_n1642) );
  OAI21_X1 Midori_rounds_U787 ( .B1(Midori_rounds_n1639), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1638), .ZN(Midori_rounds_n931)
         );
  AOI22_X1 Midori_rounds_U786 ( .A1(reset), .A2(Midori_add_Result_Start3[14]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[14]), .ZN(
        Midori_rounds_n1638) );
  XOR2_X1 Midori_rounds_U785 ( .A(Midori_rounds_SR_Inv_Result3[34]), .B(
        Midori_rounds_n1637), .Z(Midori_rounds_n1639) );
  OAI21_X1 Midori_rounds_U784 ( .B1(Midori_rounds_n1636), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1635), .ZN(
        Midori_rounds_sub_Sub_1_S2_InAff_out3[2]) );
  AOI22_X1 Midori_rounds_U783 ( .A1(reset), .A2(Midori_add_Result_Start3[15]), 
        .B1(Midori_rounds_n1255), .B2(Midori_rounds_SR_Inv_Result3[15]), .ZN(
        Midori_rounds_n1635) );
  XOR2_X1 Midori_rounds_U782 ( .A(Midori_rounds_SR_Inv_Result3[35]), .B(
        Midori_rounds_n1634), .Z(Midori_rounds_n1636) );
  OAI21_X1 Midori_rounds_U781 ( .B1(Midori_rounds_n1633), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1632), .ZN(
        Midori_rounds_sub_Sub_2_S1_InAff_out3[1]) );
  AOI22_X1 Midori_rounds_U780 ( .A1(reset), .A2(Midori_add_Result_Start3[16]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[16]), .ZN(
        Midori_rounds_n1632) );
  XOR2_X1 Midori_rounds_U779 ( .A(Midori_rounds_SR_Inv_Result3[36]), .B(
        Midori_rounds_n1631), .Z(Midori_rounds_n1633) );
  OAI21_X1 Midori_rounds_U778 ( .B1(Midori_rounds_n1630), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1629), .ZN(
        Midori_rounds_sub_Sub_2_S1_InAff_out3[0]) );
  AOI22_X1 Midori_rounds_U777 ( .A1(reset), .A2(Midori_add_Result_Start3[17]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[17]), .ZN(
        Midori_rounds_n1629) );
  XOR2_X1 Midori_rounds_U776 ( .A(Midori_rounds_SR_Inv_Result3[37]), .B(
        Midori_rounds_n1628), .Z(Midori_rounds_n1630) );
  OAI21_X1 Midori_rounds_U775 ( .B1(Midori_rounds_n1627), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1626), .ZN(Midori_rounds_n935)
         );
  AOI22_X1 Midori_rounds_U774 ( .A1(reset), .A2(Midori_add_Result_Start3[18]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[18]), .ZN(
        Midori_rounds_n1626) );
  XOR2_X1 Midori_rounds_U773 ( .A(Midori_rounds_SR_Inv_Result3[38]), .B(
        Midori_rounds_n1625), .Z(Midori_rounds_n1627) );
  OAI21_X1 Midori_rounds_U772 ( .B1(Midori_rounds_n1624), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1623), .ZN(
        Midori_rounds_sub_Sub_2_S1_InAff_out3[2]) );
  AOI22_X1 Midori_rounds_U771 ( .A1(reset), .A2(Midori_add_Result_Start3[19]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[19]), .ZN(
        Midori_rounds_n1623) );
  XOR2_X1 Midori_rounds_U770 ( .A(Midori_rounds_SR_Inv_Result3[39]), .B(
        Midori_rounds_n1622), .Z(Midori_rounds_n1624) );
  OAI21_X1 Midori_rounds_U769 ( .B1(Midori_rounds_n1621), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1620), .ZN(
        Midori_rounds_sub_Sub_2_S2_InAff_out3[1]) );
  AOI22_X1 Midori_rounds_U768 ( .A1(reset), .A2(Midori_add_Result_Start3[20]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[20]), .ZN(
        Midori_rounds_n1620) );
  XOR2_X1 Midori_rounds_U767 ( .A(Midori_rounds_SR_Inv_Result3[12]), .B(
        Midori_rounds_n1619), .Z(Midori_rounds_n1621) );
  OAI21_X1 Midori_rounds_U766 ( .B1(Midori_rounds_n1618), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1617), .ZN(
        Midori_rounds_sub_Sub_2_S2_InAff_out3[0]) );
  AOI22_X1 Midori_rounds_U765 ( .A1(reset), .A2(Midori_add_Result_Start3[21]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[21]), .ZN(
        Midori_rounds_n1617) );
  XOR2_X1 Midori_rounds_U764 ( .A(Midori_rounds_SR_Inv_Result3[13]), .B(
        Midori_rounds_n1616), .Z(Midori_rounds_n1618) );
  OAI21_X1 Midori_rounds_U763 ( .B1(Midori_rounds_n1615), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1614), .ZN(Midori_rounds_n939)
         );
  AOI22_X1 Midori_rounds_U762 ( .A1(reset), .A2(Midori_add_Result_Start3[22]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[22]), .ZN(
        Midori_rounds_n1614) );
  XOR2_X1 Midori_rounds_U761 ( .A(Midori_rounds_SR_Inv_Result3[14]), .B(
        Midori_rounds_n1613), .Z(Midori_rounds_n1615) );
  OAI21_X1 Midori_rounds_U760 ( .B1(Midori_rounds_n1612), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1611), .ZN(
        Midori_rounds_sub_Sub_2_S2_InAff_out3[2]) );
  AOI22_X1 Midori_rounds_U759 ( .A1(reset), .A2(Midori_add_Result_Start3[23]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[23]), .ZN(
        Midori_rounds_n1611) );
  XOR2_X1 Midori_rounds_U758 ( .A(Midori_rounds_SR_Inv_Result3[15]), .B(
        Midori_rounds_n1610), .Z(Midori_rounds_n1612) );
  OAI21_X1 Midori_rounds_U757 ( .B1(Midori_rounds_n1609), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1608), .ZN(
        Midori_rounds_sub_Sub_3_S1_InAff_out3[1]) );
  AOI22_X1 Midori_rounds_U756 ( .A1(reset), .A2(Midori_add_Result_Start3[24]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[24]), .ZN(
        Midori_rounds_n1608) );
  XOR2_X1 Midori_rounds_U755 ( .A(Midori_rounds_SR_Inv_Result3[48]), .B(
        Midori_rounds_n1607), .Z(Midori_rounds_n1609) );
  OAI21_X1 Midori_rounds_U754 ( .B1(Midori_rounds_n1606), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1605), .ZN(
        Midori_rounds_sub_Sub_3_S1_InAff_out3[0]) );
  AOI22_X1 Midori_rounds_U753 ( .A1(reset), .A2(Midori_add_Result_Start3[25]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[25]), .ZN(
        Midori_rounds_n1605) );
  XOR2_X1 Midori_rounds_U752 ( .A(Midori_rounds_SR_Inv_Result3[49]), .B(
        Midori_rounds_n1604), .Z(Midori_rounds_n1606) );
  OAI21_X1 Midori_rounds_U751 ( .B1(Midori_rounds_n1603), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1602), .ZN(Midori_rounds_n943)
         );
  AOI22_X1 Midori_rounds_U750 ( .A1(reset), .A2(Midori_add_Result_Start3[26]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[26]), .ZN(
        Midori_rounds_n1602) );
  XOR2_X1 Midori_rounds_U749 ( .A(Midori_rounds_SR_Inv_Result3[50]), .B(
        Midori_rounds_n1601), .Z(Midori_rounds_n1603) );
  OAI21_X1 Midori_rounds_U748 ( .B1(Midori_rounds_n1600), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1599), .ZN(
        Midori_rounds_sub_Sub_3_S1_InAff_out3[2]) );
  AOI22_X1 Midori_rounds_U747 ( .A1(reset), .A2(Midori_add_Result_Start3[27]), 
        .B1(Midori_rounds_n1254), .B2(Midori_rounds_SR_Inv_Result3[27]), .ZN(
        Midori_rounds_n1599) );
  XOR2_X1 Midori_rounds_U746 ( .A(Midori_rounds_SR_Inv_Result3[51]), .B(
        Midori_rounds_n1598), .Z(Midori_rounds_n1600) );
  OAI21_X1 Midori_rounds_U745 ( .B1(Midori_rounds_n1597), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1596), .ZN(
        Midori_rounds_sub_Sub_3_S2_InAff_out3[1]) );
  AOI22_X1 Midori_rounds_U744 ( .A1(reset), .A2(Midori_add_Result_Start3[28]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[28]), .ZN(
        Midori_rounds_n1596) );
  XOR2_X1 Midori_rounds_U743 ( .A(Midori_rounds_SR_Inv_Result3[24]), .B(
        Midori_rounds_n1595), .Z(Midori_rounds_n1597) );
  OAI21_X1 Midori_rounds_U742 ( .B1(Midori_rounds_n1594), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1593), .ZN(
        Midori_rounds_sub_Sub_3_S2_InAff_out3[0]) );
  AOI22_X1 Midori_rounds_U741 ( .A1(reset), .A2(Midori_add_Result_Start3[29]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[29]), .ZN(
        Midori_rounds_n1593) );
  XOR2_X1 Midori_rounds_U740 ( .A(Midori_rounds_SR_Inv_Result3[25]), .B(
        Midori_rounds_n1592), .Z(Midori_rounds_n1594) );
  OAI21_X1 Midori_rounds_U739 ( .B1(Midori_rounds_n1591), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1590), .ZN(Midori_rounds_n947)
         );
  AOI22_X1 Midori_rounds_U738 ( .A1(reset), .A2(Midori_add_Result_Start3[30]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[30]), .ZN(
        Midori_rounds_n1590) );
  XOR2_X1 Midori_rounds_U737 ( .A(Midori_rounds_SR_Inv_Result3[26]), .B(
        Midori_rounds_n1589), .Z(Midori_rounds_n1591) );
  OAI21_X1 Midori_rounds_U736 ( .B1(Midori_rounds_n1588), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1587), .ZN(
        Midori_rounds_sub_Sub_3_S2_InAff_out3[2]) );
  AOI22_X1 Midori_rounds_U735 ( .A1(reset), .A2(Midori_add_Result_Start3[31]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[31]), .ZN(
        Midori_rounds_n1587) );
  XOR2_X1 Midori_rounds_U734 ( .A(Midori_rounds_SR_Inv_Result3[27]), .B(
        Midori_rounds_n1586), .Z(Midori_rounds_n1588) );
  OAI21_X1 Midori_rounds_U733 ( .B1(Midori_rounds_n1585), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1584), .ZN(
        Midori_rounds_sub_Sub_4_S1_InAff_out3[1]) );
  AOI22_X1 Midori_rounds_U732 ( .A1(reset), .A2(Midori_add_Result_Start3[32]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[32]), .ZN(
        Midori_rounds_n1584) );
  XOR2_X1 Midori_rounds_U731 ( .A(Midori_rounds_SR_Inv_Result3[56]), .B(
        Midori_rounds_n1583), .Z(Midori_rounds_n1585) );
  OAI21_X1 Midori_rounds_U730 ( .B1(Midori_rounds_n1582), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1581), .ZN(
        Midori_rounds_sub_Sub_4_S1_InAff_out3[0]) );
  AOI22_X1 Midori_rounds_U729 ( .A1(reset), .A2(Midori_add_Result_Start3[33]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[33]), .ZN(
        Midori_rounds_n1581) );
  XOR2_X1 Midori_rounds_U728 ( .A(Midori_rounds_SR_Inv_Result3[57]), .B(
        Midori_rounds_n1580), .Z(Midori_rounds_n1582) );
  OAI21_X1 Midori_rounds_U727 ( .B1(Midori_rounds_n1579), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1578), .ZN(Midori_rounds_n951)
         );
  AOI22_X1 Midori_rounds_U726 ( .A1(reset), .A2(Midori_add_Result_Start3[34]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[34]), .ZN(
        Midori_rounds_n1578) );
  XOR2_X1 Midori_rounds_U725 ( .A(Midori_rounds_SR_Inv_Result3[58]), .B(
        Midori_rounds_n1577), .Z(Midori_rounds_n1579) );
  OAI21_X1 Midori_rounds_U724 ( .B1(Midori_rounds_n1576), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1575), .ZN(
        Midori_rounds_sub_Sub_4_S1_InAff_out3[2]) );
  AOI22_X1 Midori_rounds_U723 ( .A1(reset), .A2(Midori_add_Result_Start3[35]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[35]), .ZN(
        Midori_rounds_n1575) );
  XOR2_X1 Midori_rounds_U722 ( .A(Midori_rounds_SR_Inv_Result3[59]), .B(
        Midori_rounds_n1574), .Z(Midori_rounds_n1576) );
  OAI21_X1 Midori_rounds_U721 ( .B1(Midori_rounds_n1573), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1572), .ZN(
        Midori_rounds_sub_Sub_4_S2_InAff_out3[1]) );
  AOI22_X1 Midori_rounds_U720 ( .A1(reset), .A2(Midori_add_Result_Start3[36]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[36]), .ZN(
        Midori_rounds_n1572) );
  XOR2_X1 Midori_rounds_U719 ( .A(Midori_rounds_SR_Inv_Result3[16]), .B(
        Midori_rounds_n1571), .Z(Midori_rounds_n1573) );
  OAI21_X1 Midori_rounds_U718 ( .B1(Midori_rounds_n1570), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1569), .ZN(
        Midori_rounds_sub_Sub_4_S2_InAff_out3[0]) );
  AOI22_X1 Midori_rounds_U717 ( .A1(reset), .A2(Midori_add_Result_Start3[37]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[37]), .ZN(
        Midori_rounds_n1569) );
  XOR2_X1 Midori_rounds_U716 ( .A(Midori_rounds_SR_Inv_Result3[17]), .B(
        Midori_rounds_n1568), .Z(Midori_rounds_n1570) );
  OAI21_X1 Midori_rounds_U715 ( .B1(Midori_rounds_n1567), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1566), .ZN(Midori_rounds_n955)
         );
  AOI22_X1 Midori_rounds_U714 ( .A1(reset), .A2(Midori_add_Result_Start3[38]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[38]), .ZN(
        Midori_rounds_n1566) );
  XOR2_X1 Midori_rounds_U713 ( .A(Midori_rounds_SR_Inv_Result3[18]), .B(
        Midori_rounds_n1565), .Z(Midori_rounds_n1567) );
  OAI21_X1 Midori_rounds_U712 ( .B1(Midori_rounds_n1564), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1563), .ZN(
        Midori_rounds_sub_Sub_4_S2_InAff_out3[2]) );
  AOI22_X1 Midori_rounds_U711 ( .A1(reset), .A2(Midori_add_Result_Start3[39]), 
        .B1(Midori_rounds_n1253), .B2(Midori_rounds_SR_Inv_Result3[39]), .ZN(
        Midori_rounds_n1563) );
  XOR2_X1 Midori_rounds_U710 ( .A(Midori_rounds_SR_Inv_Result3[19]), .B(
        Midori_rounds_n1562), .Z(Midori_rounds_n1564) );
  OAI21_X1 Midori_rounds_U709 ( .B1(Midori_rounds_n1561), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1560), .ZN(
        Midori_rounds_sub_Sub_5_S1_InAff_out3[1]) );
  AOI22_X1 Midori_rounds_U708 ( .A1(reset), .A2(Midori_add_Result_Start3[40]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[40]), .ZN(
        Midori_rounds_n1560) );
  XOR2_X1 Midori_rounds_U707 ( .A(Midori_rounds_SR_Inv_Result3[44]), .B(
        Midori_rounds_n1559), .Z(Midori_rounds_n1561) );
  OAI21_X1 Midori_rounds_U706 ( .B1(Midori_rounds_n1558), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1557), .ZN(
        Midori_rounds_sub_Sub_5_S1_InAff_out3[0]) );
  AOI22_X1 Midori_rounds_U705 ( .A1(reset), .A2(Midori_add_Result_Start3[41]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[41]), .ZN(
        Midori_rounds_n1557) );
  XOR2_X1 Midori_rounds_U704 ( .A(Midori_rounds_SR_Inv_Result3[45]), .B(
        Midori_rounds_n1556), .Z(Midori_rounds_n1558) );
  OAI21_X1 Midori_rounds_U703 ( .B1(Midori_rounds_n1555), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1554), .ZN(Midori_rounds_n959)
         );
  AOI22_X1 Midori_rounds_U702 ( .A1(reset), .A2(Midori_add_Result_Start3[42]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[42]), .ZN(
        Midori_rounds_n1554) );
  XOR2_X1 Midori_rounds_U701 ( .A(Midori_rounds_SR_Inv_Result3[46]), .B(
        Midori_rounds_n1553), .Z(Midori_rounds_n1555) );
  OAI21_X1 Midori_rounds_U700 ( .B1(Midori_rounds_n1552), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1551), .ZN(
        Midori_rounds_sub_Sub_5_S1_InAff_out3[2]) );
  AOI22_X1 Midori_rounds_U699 ( .A1(reset), .A2(Midori_add_Result_Start3[43]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[43]), .ZN(
        Midori_rounds_n1551) );
  XOR2_X1 Midori_rounds_U698 ( .A(Midori_rounds_SR_Inv_Result3[47]), .B(
        Midori_rounds_n1550), .Z(Midori_rounds_n1552) );
  OAI21_X1 Midori_rounds_U697 ( .B1(Midori_rounds_n1549), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1548), .ZN(
        Midori_rounds_sub_Sub_5_S2_InAff_out3[1]) );
  AOI22_X1 Midori_rounds_U696 ( .A1(reset), .A2(Midori_add_Result_Start3[44]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[44]), .ZN(
        Midori_rounds_n1548) );
  XOR2_X1 Midori_rounds_U695 ( .A(Midori_rounds_SR_Inv_Result3[4]), .B(
        Midori_rounds_n1547), .Z(Midori_rounds_n1549) );
  OAI21_X1 Midori_rounds_U694 ( .B1(Midori_rounds_n1546), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1545), .ZN(
        Midori_rounds_sub_Sub_5_S2_InAff_out3[0]) );
  AOI22_X1 Midori_rounds_U693 ( .A1(reset), .A2(Midori_add_Result_Start3[45]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[45]), .ZN(
        Midori_rounds_n1545) );
  XOR2_X1 Midori_rounds_U692 ( .A(Midori_rounds_SR_Inv_Result3[5]), .B(
        Midori_rounds_n1544), .Z(Midori_rounds_n1546) );
  OAI21_X1 Midori_rounds_U691 ( .B1(Midori_rounds_n1543), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1542), .ZN(Midori_rounds_n963)
         );
  AOI22_X1 Midori_rounds_U690 ( .A1(reset), .A2(Midori_add_Result_Start3[46]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[46]), .ZN(
        Midori_rounds_n1542) );
  XOR2_X1 Midori_rounds_U689 ( .A(Midori_rounds_SR_Inv_Result3[6]), .B(
        Midori_rounds_n1541), .Z(Midori_rounds_n1543) );
  OAI21_X1 Midori_rounds_U688 ( .B1(Midori_rounds_n1540), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1539), .ZN(
        Midori_rounds_sub_Sub_5_S2_InAff_out3[2]) );
  AOI22_X1 Midori_rounds_U687 ( .A1(reset), .A2(Midori_add_Result_Start3[47]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[47]), .ZN(
        Midori_rounds_n1539) );
  XOR2_X1 Midori_rounds_U686 ( .A(Midori_rounds_SR_Inv_Result3[7]), .B(
        Midori_rounds_n1538), .Z(Midori_rounds_n1540) );
  OAI21_X1 Midori_rounds_U685 ( .B1(Midori_rounds_n1537), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1536), .ZN(
        Midori_rounds_sub_Sub_6_S1_InAff_out3[1]) );
  AOI22_X1 Midori_rounds_U684 ( .A1(reset), .A2(Midori_add_Result_Start3[48]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[48]), .ZN(
        Midori_rounds_n1536) );
  XOR2_X1 Midori_rounds_U683 ( .A(Midori_rounds_SR_Inv_Result3[0]), .B(
        Midori_rounds_n1535), .Z(Midori_rounds_n1537) );
  OAI21_X1 Midori_rounds_U682 ( .B1(Midori_rounds_n1534), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1533), .ZN(
        Midori_rounds_sub_Sub_6_S1_InAff_out3[0]) );
  AOI22_X1 Midori_rounds_U681 ( .A1(reset), .A2(Midori_add_Result_Start3[49]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[49]), .ZN(
        Midori_rounds_n1533) );
  XOR2_X1 Midori_rounds_U680 ( .A(Midori_rounds_SR_Inv_Result3[1]), .B(
        Midori_rounds_n1532), .Z(Midori_rounds_n1534) );
  OAI21_X1 Midori_rounds_U679 ( .B1(Midori_rounds_n1531), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1530), .ZN(Midori_rounds_n967)
         );
  AOI22_X1 Midori_rounds_U678 ( .A1(reset), .A2(Midori_add_Result_Start3[50]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[50]), .ZN(
        Midori_rounds_n1530) );
  XOR2_X1 Midori_rounds_U677 ( .A(Midori_rounds_SR_Inv_Result3[2]), .B(
        Midori_rounds_n1529), .Z(Midori_rounds_n1531) );
  OAI21_X1 Midori_rounds_U676 ( .B1(Midori_rounds_n1528), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1527), .ZN(
        Midori_rounds_sub_Sub_6_S1_InAff_out3[2]) );
  AOI22_X1 Midori_rounds_U675 ( .A1(reset), .A2(Midori_add_Result_Start3[51]), 
        .B1(Midori_rounds_n1252), .B2(Midori_rounds_SR_Inv_Result3[51]), .ZN(
        Midori_rounds_n1527) );
  XOR2_X1 Midori_rounds_U674 ( .A(Midori_rounds_SR_Inv_Result3[3]), .B(
        Midori_rounds_n1526), .Z(Midori_rounds_n1528) );
  OAI21_X1 Midori_rounds_U673 ( .B1(Midori_rounds_n1525), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1524), .ZN(
        Midori_rounds_sub_Sub_6_S2_InAff_out3[1]) );
  AOI22_X1 Midori_rounds_U672 ( .A1(reset), .A2(Midori_add_Result_Start3[52]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[52]), .ZN(
        Midori_rounds_n1524) );
  XOR2_X1 Midori_rounds_U671 ( .A(Midori_rounds_SR_Inv_Result3[40]), .B(
        Midori_rounds_n1523), .Z(Midori_rounds_n1525) );
  OAI21_X1 Midori_rounds_U670 ( .B1(Midori_rounds_n1522), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1521), .ZN(
        Midori_rounds_sub_Sub_6_S2_InAff_out3[0]) );
  AOI22_X1 Midori_rounds_U669 ( .A1(reset), .A2(Midori_add_Result_Start3[53]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[53]), .ZN(
        Midori_rounds_n1521) );
  XOR2_X1 Midori_rounds_U668 ( .A(Midori_rounds_SR_Inv_Result3[41]), .B(
        Midori_rounds_n1520), .Z(Midori_rounds_n1522) );
  OAI21_X1 Midori_rounds_U667 ( .B1(Midori_rounds_n1519), .B2(
        Midori_rounds_n1262), .A(Midori_rounds_n1518), .ZN(Midori_rounds_n971)
         );
  AOI22_X1 Midori_rounds_U666 ( .A1(reset), .A2(Midori_add_Result_Start3[54]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[54]), .ZN(
        Midori_rounds_n1518) );
  XOR2_X1 Midori_rounds_U665 ( .A(Midori_rounds_SR_Inv_Result3[42]), .B(
        Midori_rounds_n1517), .Z(Midori_rounds_n1519) );
  OAI21_X1 Midori_rounds_U664 ( .B1(Midori_rounds_n1516), .B2(
        Midori_rounds_n1263), .A(Midori_rounds_n1515), .ZN(
        Midori_rounds_sub_Sub_6_S2_InAff_out3[2]) );
  AOI22_X1 Midori_rounds_U663 ( .A1(reset), .A2(Midori_add_Result_Start3[55]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[55]), .ZN(
        Midori_rounds_n1515) );
  XOR2_X1 Midori_rounds_U662 ( .A(Midori_rounds_SR_Inv_Result3[43]), .B(
        Midori_rounds_n1514), .Z(Midori_rounds_n1516) );
  OAI21_X1 Midori_rounds_U661 ( .B1(Midori_rounds_n1513), .B2(
        Midori_rounds_n1264), .A(Midori_rounds_n1512), .ZN(
        Midori_rounds_sub_Sub_7_S1_InAff_out3[1]) );
  AOI22_X1 Midori_rounds_U660 ( .A1(reset), .A2(Midori_add_Result_Start3[56]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[56]), .ZN(
        Midori_rounds_n1512) );
  XOR2_X1 Midori_rounds_U659 ( .A(Midori_rounds_SR_Inv_Result3[20]), .B(
        Midori_rounds_n1511), .Z(Midori_rounds_n1513) );
  OAI21_X1 Midori_rounds_U658 ( .B1(Midori_rounds_n1510), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1509), .ZN(
        Midori_rounds_sub_Sub_7_S1_InAff_out3[0]) );
  AOI22_X1 Midori_rounds_U657 ( .A1(reset), .A2(Midori_add_Result_Start3[57]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[57]), .ZN(
        Midori_rounds_n1509) );
  XOR2_X1 Midori_rounds_U656 ( .A(Midori_rounds_SR_Inv_Result3[21]), .B(
        Midori_rounds_n1508), .Z(Midori_rounds_n1510) );
  OAI21_X1 Midori_rounds_U655 ( .B1(Midori_rounds_n1507), .B2(
        Midori_rounds_n1261), .A(Midori_rounds_n1506), .ZN(Midori_rounds_n975)
         );
  AOI22_X1 Midori_rounds_U654 ( .A1(reset), .A2(Midori_add_Result_Start3[58]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[58]), .ZN(
        Midori_rounds_n1506) );
  XOR2_X1 Midori_rounds_U653 ( .A(Midori_rounds_SR_Inv_Result3[22]), .B(
        Midori_rounds_n1505), .Z(Midori_rounds_n1507) );
  OAI21_X1 Midori_rounds_U652 ( .B1(Midori_rounds_n1504), .B2(
        Midori_rounds_n1260), .A(Midori_rounds_n1503), .ZN(
        Midori_rounds_sub_Sub_7_S1_InAff_out3[2]) );
  AOI22_X1 Midori_rounds_U651 ( .A1(reset), .A2(Midori_add_Result_Start3[59]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[59]), .ZN(
        Midori_rounds_n1503) );
  XOR2_X1 Midori_rounds_U650 ( .A(Midori_rounds_SR_Inv_Result3[23]), .B(
        Midori_rounds_n1502), .Z(Midori_rounds_n1504) );
  OAI21_X1 Midori_rounds_U649 ( .B1(Midori_rounds_n1501), .B2(
        Midori_rounds_n1266), .A(Midori_rounds_n1500), .ZN(
        Midori_rounds_sub_Sub_7_S2_InAff_out3[1]) );
  AOI22_X1 Midori_rounds_U648 ( .A1(reset), .A2(Midori_add_Result_Start3[60]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[60]), .ZN(
        Midori_rounds_n1500) );
  XOR2_X1 Midori_rounds_U647 ( .A(Midori_rounds_SR_Inv_Result3[60]), .B(
        Midori_rounds_n1499), .Z(Midori_rounds_n1501) );
  OAI21_X1 Midori_rounds_U646 ( .B1(Midori_rounds_n1498), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1497), .ZN(
        Midori_rounds_sub_Sub_7_S2_InAff_out3[0]) );
  AOI22_X1 Midori_rounds_U645 ( .A1(reset), .A2(Midori_add_Result_Start3[61]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[61]), .ZN(
        Midori_rounds_n1497) );
  XOR2_X1 Midori_rounds_U644 ( .A(Midori_rounds_SR_Inv_Result3[61]), .B(
        Midori_rounds_n1496), .Z(Midori_rounds_n1498) );
  OAI21_X1 Midori_rounds_U643 ( .B1(Midori_rounds_n1495), .B2(
        Midori_rounds_n2066), .A(Midori_rounds_n1494), .ZN(Midori_rounds_n979)
         );
  AOI22_X1 Midori_rounds_U642 ( .A1(reset), .A2(Midori_add_Result_Start3[62]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[62]), .ZN(
        Midori_rounds_n1494) );
  XOR2_X1 Midori_rounds_U641 ( .A(Midori_rounds_SR_Inv_Result3[62]), .B(
        Midori_rounds_n1493), .Z(Midori_rounds_n1495) );
  OAI21_X1 Midori_rounds_U640 ( .B1(Midori_rounds_n1492), .B2(
        Midori_rounds_n1265), .A(Midori_rounds_n1491), .ZN(
        Midori_rounds_sub_Sub_7_S2_InAff_out3[2]) );
  AOI22_X1 Midori_rounds_U639 ( .A1(reset), .A2(Midori_add_Result_Start3[63]), 
        .B1(Midori_rounds_n1251), .B2(Midori_rounds_SR_Inv_Result3[63]), .ZN(
        Midori_rounds_n1491) );
  XOR2_X1 Midori_rounds_U638 ( .A(Midori_rounds_SR_Inv_Result3[63]), .B(
        Midori_rounds_n1489), .Z(Midori_rounds_n1492) );
  MUX2_X1 Midori_rounds_U637 ( .A(Midori_rounds_n1488), .B(
        Midori_rounds_SR_Result3[9]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[9]) );
  XNOR2_X1 Midori_rounds_U636 ( .A(Midori_rounds_SR_Result3[9]), .B(
        Midori_rounds_n1652), .ZN(Midori_rounds_n1488) );
  AOI22_X1 Midori_rounds_U635 ( .A1(Midori_rounds_n1270), .A2(Key3[9]), .B1(
        Key3[73]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1652) );
  MUX2_X1 Midori_rounds_U634 ( .A(Midori_rounds_n1487), .B(
        Midori_rounds_SR_Result3[8]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[8]) );
  XNOR2_X1 Midori_rounds_U633 ( .A(Midori_rounds_SR_Result3[8]), .B(
        Midori_rounds_n1655), .ZN(Midori_rounds_n1487) );
  AOI22_X1 Midori_rounds_U632 ( .A1(Midori_rounds_n1270), .A2(Key3[8]), .B1(
        Key3[72]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1655) );
  MUX2_X1 Midori_rounds_U631 ( .A(Midori_rounds_n1486), .B(
        Midori_rounds_SR_Result3[7]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[7]) );
  XNOR2_X1 Midori_rounds_U630 ( .A(Midori_rounds_SR_Result3[47]), .B(
        Midori_rounds_n1658), .ZN(Midori_rounds_n1486) );
  AOI22_X1 Midori_rounds_U629 ( .A1(Midori_rounds_n1268), .A2(Key3[7]), .B1(
        Key3[71]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1658) );
  MUX2_X1 Midori_rounds_U628 ( .A(Midori_rounds_n1485), .B(
        Midori_rounds_SR_Result3[6]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[6]) );
  XNOR2_X1 Midori_rounds_U627 ( .A(Midori_rounds_SR_Result3[46]), .B(
        Midori_rounds_n1661), .ZN(Midori_rounds_n1485) );
  AOI22_X1 Midori_rounds_U626 ( .A1(Midori_rounds_n1273), .A2(Key3[6]), .B1(
        Key3[70]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1661) );
  MUX2_X1 Midori_rounds_U625 ( .A(Midori_rounds_n1484), .B(
        Midori_rounds_SR_Result3[63]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[63]) );
  XNOR2_X1 Midori_rounds_U624 ( .A(Midori_rounds_SR_Result3[63]), .B(
        Midori_rounds_n1489), .ZN(Midori_rounds_n1484) );
  AOI22_X1 Midori_rounds_U623 ( .A1(Midori_rounds_n1271), .A2(Key3[63]), .B1(
        Key3[127]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1489) );
  MUX2_X1 Midori_rounds_U622 ( .A(Midori_rounds_n1483), .B(
        Midori_rounds_SR_Result3[62]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[62]) );
  XNOR2_X1 Midori_rounds_U621 ( .A(Midori_rounds_SR_Result3[62]), .B(
        Midori_rounds_n1493), .ZN(Midori_rounds_n1483) );
  AOI22_X1 Midori_rounds_U620 ( .A1(Midori_rounds_n1274), .A2(Key3[62]), .B1(
        Key3[126]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1493) );
  MUX2_X1 Midori_rounds_U619 ( .A(Midori_rounds_n1482), .B(
        Midori_rounds_SR_Result3[61]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[61]) );
  XNOR2_X1 Midori_rounds_U618 ( .A(Midori_rounds_SR_Result3[61]), .B(
        Midori_rounds_n1496), .ZN(Midori_rounds_n1482) );
  AOI22_X1 Midori_rounds_U617 ( .A1(Midori_rounds_n1272), .A2(Key3[61]), .B1(
        Key3[125]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1496) );
  MUX2_X1 Midori_rounds_U616 ( .A(Midori_rounds_n1481), .B(
        Midori_rounds_SR_Result3[60]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[60]) );
  XNOR2_X1 Midori_rounds_U615 ( .A(Midori_rounds_SR_Result3[60]), .B(
        Midori_rounds_n1499), .ZN(Midori_rounds_n1481) );
  AOI22_X1 Midori_rounds_U614 ( .A1(Midori_rounds_n1271), .A2(Key3[60]), .B1(
        Key3[124]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1499) );
  MUX2_X1 Midori_rounds_U613 ( .A(Midori_rounds_n1480), .B(
        Midori_rounds_SR_Result3[5]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[5]) );
  XNOR2_X1 Midori_rounds_U612 ( .A(Midori_rounds_SR_Result3[45]), .B(
        Midori_rounds_n1664), .ZN(Midori_rounds_n1480) );
  AOI22_X1 Midori_rounds_U611 ( .A1(Midori_rounds_n1271), .A2(Key3[5]), .B1(
        Key3[69]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1664) );
  MUX2_X1 Midori_rounds_U610 ( .A(Midori_rounds_n1479), .B(
        Midori_rounds_SR_Result3[59]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[59]) );
  XNOR2_X1 Midori_rounds_U609 ( .A(Midori_rounds_SR_Result3[35]), .B(
        Midori_rounds_n1502), .ZN(Midori_rounds_n1479) );
  AOI22_X1 Midori_rounds_U608 ( .A1(Midori_rounds_n1269), .A2(Key3[59]), .B1(
        Key3[123]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1502) );
  MUX2_X1 Midori_rounds_U607 ( .A(Midori_rounds_n1478), .B(
        Midori_rounds_SR_Result3[58]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[58]) );
  XNOR2_X1 Midori_rounds_U606 ( .A(Midori_rounds_SR_Result3[34]), .B(
        Midori_rounds_n1505), .ZN(Midori_rounds_n1478) );
  AOI22_X1 Midori_rounds_U605 ( .A1(Midori_rounds_n1272), .A2(Key3[58]), .B1(
        Key3[122]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1505) );
  MUX2_X1 Midori_rounds_U604 ( .A(Midori_rounds_n1477), .B(
        Midori_rounds_SR_Result3[57]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[57]) );
  XNOR2_X1 Midori_rounds_U603 ( .A(Midori_rounds_SR_Result3[33]), .B(
        Midori_rounds_n1508), .ZN(Midori_rounds_n1477) );
  AOI22_X1 Midori_rounds_U602 ( .A1(Midori_rounds_n1274), .A2(Key3[57]), .B1(
        Key3[121]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1508) );
  MUX2_X1 Midori_rounds_U601 ( .A(Midori_rounds_n1476), .B(
        Midori_rounds_SR_Result3[56]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input3[56]) );
  XNOR2_X1 Midori_rounds_U600 ( .A(Midori_rounds_SR_Result3[32]), .B(
        Midori_rounds_n1511), .ZN(Midori_rounds_n1476) );
  AOI22_X1 Midori_rounds_U599 ( .A1(Midori_rounds_n1271), .A2(Key3[56]), .B1(
        Key3[120]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1511) );
  MUX2_X1 Midori_rounds_U598 ( .A(Midori_rounds_n1475), .B(
        Midori_rounds_SR_Result3[55]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input3[55]) );
  XNOR2_X1 Midori_rounds_U597 ( .A(Midori_rounds_SR_Result3[7]), .B(
        Midori_rounds_n1514), .ZN(Midori_rounds_n1475) );
  AOI22_X1 Midori_rounds_U596 ( .A1(Midori_rounds_n1270), .A2(Key3[55]), .B1(
        Key3[119]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1514) );
  MUX2_X1 Midori_rounds_U595 ( .A(Midori_rounds_n1474), .B(
        Midori_rounds_SR_Result3[54]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[54]) );
  XNOR2_X1 Midori_rounds_U594 ( .A(Midori_rounds_SR_Result3[6]), .B(
        Midori_rounds_n1517), .ZN(Midori_rounds_n1474) );
  AOI22_X1 Midori_rounds_U593 ( .A1(Midori_rounds_n1274), .A2(Key3[54]), .B1(
        Key3[118]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1517) );
  MUX2_X1 Midori_rounds_U592 ( .A(Midori_rounds_n1473), .B(
        Midori_rounds_SR_Result3[53]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input3[53]) );
  XNOR2_X1 Midori_rounds_U591 ( .A(Midori_rounds_SR_Result3[5]), .B(
        Midori_rounds_n1520), .ZN(Midori_rounds_n1473) );
  AOI22_X1 Midori_rounds_U590 ( .A1(Midori_rounds_n1270), .A2(Key3[53]), .B1(
        Key3[117]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1520) );
  MUX2_X1 Midori_rounds_U589 ( .A(Midori_rounds_n1472), .B(
        Midori_rounds_SR_Result3[52]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input3[52]) );
  XNOR2_X1 Midori_rounds_U588 ( .A(Midori_rounds_SR_Result3[4]), .B(
        Midori_rounds_n1523), .ZN(Midori_rounds_n1472) );
  AOI22_X1 Midori_rounds_U587 ( .A1(Midori_rounds_n1272), .A2(Key3[52]), .B1(
        Key3[116]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1523) );
  MUX2_X1 Midori_rounds_U586 ( .A(Midori_rounds_n1471), .B(
        Midori_rounds_SR_Result3[51]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input3[51]) );
  XNOR2_X1 Midori_rounds_U585 ( .A(Midori_rounds_SR_Result3[27]), .B(
        Midori_rounds_n1526), .ZN(Midori_rounds_n1471) );
  AOI22_X1 Midori_rounds_U584 ( .A1(Midori_rounds_n1272), .A2(Key3[51]), .B1(
        Key3[115]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1526) );
  MUX2_X1 Midori_rounds_U583 ( .A(Midori_rounds_n1470), .B(
        Midori_rounds_SR_Result3[50]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input3[50]) );
  XNOR2_X1 Midori_rounds_U582 ( .A(Midori_rounds_SR_Result3[26]), .B(
        Midori_rounds_n1529), .ZN(Midori_rounds_n1470) );
  AOI22_X1 Midori_rounds_U581 ( .A1(Midori_rounds_n1268), .A2(Key3[50]), .B1(
        Key3[114]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1529) );
  MUX2_X1 Midori_rounds_U580 ( .A(Midori_rounds_n1469), .B(
        Midori_rounds_SR_Result3[4]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[4]) );
  XNOR2_X1 Midori_rounds_U579 ( .A(Midori_rounds_SR_Result3[44]), .B(
        Midori_rounds_n1667), .ZN(Midori_rounds_n1469) );
  AOI22_X1 Midori_rounds_U578 ( .A1(Midori_rounds_n1273), .A2(Key3[4]), .B1(
        Key3[68]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1667) );
  MUX2_X1 Midori_rounds_U577 ( .A(Midori_rounds_n1468), .B(
        Midori_rounds_SR_Result3[49]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[49]) );
  XNOR2_X1 Midori_rounds_U576 ( .A(Midori_rounds_SR_Result3[25]), .B(
        Midori_rounds_n1532), .ZN(Midori_rounds_n1468) );
  AOI22_X1 Midori_rounds_U575 ( .A1(Midori_rounds_n1268), .A2(Key3[49]), .B1(
        Key3[113]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1532) );
  MUX2_X1 Midori_rounds_U574 ( .A(Midori_rounds_n1467), .B(
        Midori_rounds_SR_Result3[48]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input3[48]) );
  XNOR2_X1 Midori_rounds_U573 ( .A(Midori_rounds_SR_Result3[24]), .B(
        Midori_rounds_n1535), .ZN(Midori_rounds_n1467) );
  AOI22_X1 Midori_rounds_U572 ( .A1(Midori_rounds_n1272), .A2(Key3[48]), .B1(
        Key3[112]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1535) );
  MUX2_X1 Midori_rounds_U571 ( .A(Midori_rounds_n1466), .B(
        Midori_rounds_SR_Result3[47]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input3[47]) );
  XNOR2_X1 Midori_rounds_U570 ( .A(Midori_rounds_SR_Result3[43]), .B(
        Midori_rounds_n1538), .ZN(Midori_rounds_n1466) );
  AOI22_X1 Midori_rounds_U569 ( .A1(Midori_rounds_n1273), .A2(Key3[47]), .B1(
        Key3[111]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1538) );
  MUX2_X1 Midori_rounds_U568 ( .A(Midori_rounds_n1465), .B(
        Midori_rounds_SR_Result3[46]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input3[46]) );
  XNOR2_X1 Midori_rounds_U567 ( .A(Midori_rounds_SR_Result3[42]), .B(
        Midori_rounds_n1541), .ZN(Midori_rounds_n1465) );
  AOI22_X1 Midori_rounds_U566 ( .A1(Midori_rounds_n1268), .A2(Key3[46]), .B1(
        Key3[110]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1541) );
  MUX2_X1 Midori_rounds_U565 ( .A(Midori_rounds_n1464), .B(
        Midori_rounds_SR_Result3[45]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[45]) );
  XNOR2_X1 Midori_rounds_U564 ( .A(Midori_rounds_SR_Result3[41]), .B(
        Midori_rounds_n1544), .ZN(Midori_rounds_n1464) );
  AOI22_X1 Midori_rounds_U563 ( .A1(Midori_rounds_n1269), .A2(Key3[45]), .B1(
        Key3[109]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1544) );
  MUX2_X1 Midori_rounds_U562 ( .A(Midori_rounds_n1463), .B(
        Midori_rounds_SR_Result3[44]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input3[44]) );
  XNOR2_X1 Midori_rounds_U561 ( .A(Midori_rounds_SR_Result3[40]), .B(
        Midori_rounds_n1547), .ZN(Midori_rounds_n1463) );
  AOI22_X1 Midori_rounds_U560 ( .A1(Midori_rounds_n1274), .A2(Key3[44]), .B1(
        Key3[108]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1547) );
  MUX2_X1 Midori_rounds_U559 ( .A(Midori_rounds_n1462), .B(
        Midori_rounds_SR_Result3[43]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[43]) );
  XNOR2_X1 Midori_rounds_U558 ( .A(Midori_rounds_SR_Result3[55]), .B(
        Midori_rounds_n1550), .ZN(Midori_rounds_n1462) );
  AOI22_X1 Midori_rounds_U557 ( .A1(Midori_rounds_n1269), .A2(Key3[43]), .B1(
        Key3[107]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1550) );
  MUX2_X1 Midori_rounds_U556 ( .A(Midori_rounds_n1461), .B(
        Midori_rounds_SR_Result3[42]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input3[42]) );
  XNOR2_X1 Midori_rounds_U555 ( .A(Midori_rounds_SR_Result3[54]), .B(
        Midori_rounds_n1553), .ZN(Midori_rounds_n1461) );
  AOI22_X1 Midori_rounds_U554 ( .A1(Midori_rounds_n1269), .A2(Key3[42]), .B1(
        Key3[106]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1553) );
  MUX2_X1 Midori_rounds_U553 ( .A(Midori_rounds_n1460), .B(
        Midori_rounds_SR_Result3[41]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[41]) );
  XNOR2_X1 Midori_rounds_U552 ( .A(Midori_rounds_SR_Result3[53]), .B(
        Midori_rounds_n1556), .ZN(Midori_rounds_n1460) );
  AOI22_X1 Midori_rounds_U551 ( .A1(Midori_rounds_n1269), .A2(Key3[41]), .B1(
        Key3[105]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1556) );
  MUX2_X1 Midori_rounds_U550 ( .A(Midori_rounds_n1459), .B(
        Midori_rounds_SR_Result3[40]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[40]) );
  XNOR2_X1 Midori_rounds_U549 ( .A(Midori_rounds_SR_Result3[52]), .B(
        Midori_rounds_n1559), .ZN(Midori_rounds_n1459) );
  AOI22_X1 Midori_rounds_U548 ( .A1(Midori_rounds_n1272), .A2(Key3[40]), .B1(
        Key3[104]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1559) );
  MUX2_X1 Midori_rounds_U547 ( .A(Midori_rounds_n1458), .B(
        Midori_rounds_SR_Result3[3]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input3[3]) );
  XNOR2_X1 Midori_rounds_U546 ( .A(Midori_rounds_SR_Result3[51]), .B(
        Midori_rounds_n1670), .ZN(Midori_rounds_n1458) );
  AOI22_X1 Midori_rounds_U545 ( .A1(Midori_rounds_n1269), .A2(Key3[3]), .B1(
        Key3[67]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1670) );
  MUX2_X1 Midori_rounds_U544 ( .A(Midori_rounds_n1457), .B(
        Midori_rounds_SR_Result3[39]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[39]) );
  XNOR2_X1 Midori_rounds_U543 ( .A(Midori_rounds_SR_Result3[19]), .B(
        Midori_rounds_n1562), .ZN(Midori_rounds_n1457) );
  AOI22_X1 Midori_rounds_U542 ( .A1(Midori_rounds_n1268), .A2(Key3[39]), .B1(
        Key3[103]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1562) );
  MUX2_X1 Midori_rounds_U541 ( .A(Midori_rounds_n1456), .B(
        Midori_rounds_SR_Result3[38]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[38]) );
  XNOR2_X1 Midori_rounds_U540 ( .A(Midori_rounds_SR_Result3[18]), .B(
        Midori_rounds_n1565), .ZN(Midori_rounds_n1456) );
  AOI22_X1 Midori_rounds_U539 ( .A1(Midori_rounds_n1268), .A2(Key3[38]), .B1(
        Key3[102]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1565) );
  MUX2_X1 Midori_rounds_U538 ( .A(Midori_rounds_n1455), .B(
        Midori_rounds_SR_Result3[37]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[37]) );
  XNOR2_X1 Midori_rounds_U537 ( .A(Midori_rounds_SR_Result3[17]), .B(
        Midori_rounds_n1568), .ZN(Midori_rounds_n1455) );
  AOI22_X1 Midori_rounds_U536 ( .A1(Midori_rounds_n1268), .A2(Key3[37]), .B1(
        Key3[101]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1568) );
  MUX2_X1 Midori_rounds_U535 ( .A(Midori_rounds_n1454), .B(
        Midori_rounds_SR_Result3[36]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input3[36]) );
  XNOR2_X1 Midori_rounds_U534 ( .A(Midori_rounds_SR_Result3[16]), .B(
        Midori_rounds_n1571), .ZN(Midori_rounds_n1454) );
  AOI22_X1 Midori_rounds_U533 ( .A1(Midori_rounds_n1273), .A2(Key3[36]), .B1(
        Key3[100]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1571) );
  MUX2_X1 Midori_rounds_U532 ( .A(Midori_rounds_n1453), .B(
        Midori_rounds_SR_Result3[35]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[35]) );
  XNOR2_X1 Midori_rounds_U531 ( .A(Midori_rounds_SR_Result3[15]), .B(
        Midori_rounds_n1574), .ZN(Midori_rounds_n1453) );
  AOI22_X1 Midori_rounds_U530 ( .A1(Midori_rounds_n1268), .A2(Key3[35]), .B1(
        Key3[99]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1574) );
  MUX2_X1 Midori_rounds_U529 ( .A(Midori_rounds_n1452), .B(
        Midori_rounds_SR_Result3[34]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input3[34]) );
  XNOR2_X1 Midori_rounds_U528 ( .A(Midori_rounds_SR_Result3[14]), .B(
        Midori_rounds_n1577), .ZN(Midori_rounds_n1452) );
  AOI22_X1 Midori_rounds_U527 ( .A1(Midori_rounds_n1269), .A2(Key3[34]), .B1(
        Key3[98]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1577) );
  MUX2_X1 Midori_rounds_U526 ( .A(Midori_rounds_n1451), .B(
        Midori_rounds_SR_Result3[33]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input3[33]) );
  XNOR2_X1 Midori_rounds_U525 ( .A(Midori_rounds_SR_Result3[13]), .B(
        Midori_rounds_n1580), .ZN(Midori_rounds_n1451) );
  AOI22_X1 Midori_rounds_U524 ( .A1(Midori_rounds_n1274), .A2(Key3[33]), .B1(
        Key3[97]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1580) );
  MUX2_X1 Midori_rounds_U523 ( .A(Midori_rounds_n1450), .B(
        Midori_rounds_SR_Result3[32]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input3[32]) );
  XNOR2_X1 Midori_rounds_U522 ( .A(Midori_rounds_SR_Result3[12]), .B(
        Midori_rounds_n1583), .ZN(Midori_rounds_n1450) );
  AOI22_X1 Midori_rounds_U521 ( .A1(Midori_rounds_n1274), .A2(Key3[32]), .B1(
        Key3[96]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1583) );
  MUX2_X1 Midori_rounds_U520 ( .A(Midori_rounds_n1449), .B(
        Midori_rounds_SR_Result3[31]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[31]) );
  XNOR2_X1 Midori_rounds_U519 ( .A(Midori_rounds_SR_Result3[3]), .B(
        Midori_rounds_n1586), .ZN(Midori_rounds_n1449) );
  AOI22_X1 Midori_rounds_U518 ( .A1(Midori_rounds_n1274), .A2(Key3[31]), .B1(
        Key3[95]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1586) );
  MUX2_X1 Midori_rounds_U517 ( .A(Midori_rounds_n1448), .B(
        Midori_rounds_SR_Result3[30]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input3[30]) );
  XNOR2_X1 Midori_rounds_U516 ( .A(Midori_rounds_SR_Result3[2]), .B(
        Midori_rounds_n1589), .ZN(Midori_rounds_n1448) );
  AOI22_X1 Midori_rounds_U515 ( .A1(Midori_rounds_n1274), .A2(Key3[30]), .B1(
        Key3[94]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1589) );
  MUX2_X1 Midori_rounds_U514 ( .A(Midori_rounds_n1447), .B(
        Midori_rounds_SR_Result3[2]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input3[2]) );
  XNOR2_X1 Midori_rounds_U513 ( .A(Midori_rounds_SR_Result3[50]), .B(
        Midori_rounds_n1673), .ZN(Midori_rounds_n1447) );
  AOI22_X1 Midori_rounds_U512 ( .A1(Midori_rounds_n1274), .A2(Key3[2]), .B1(
        Key3[66]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1673) );
  MUX2_X1 Midori_rounds_U511 ( .A(Midori_rounds_n1446), .B(
        Midori_rounds_SR_Result3[29]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[29]) );
  XNOR2_X1 Midori_rounds_U510 ( .A(Midori_rounds_SR_Result3[1]), .B(
        Midori_rounds_n1592), .ZN(Midori_rounds_n1446) );
  AOI22_X1 Midori_rounds_U509 ( .A1(Midori_rounds_n1274), .A2(Key3[29]), .B1(
        Key3[93]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1592) );
  MUX2_X1 Midori_rounds_U508 ( .A(Midori_rounds_n1445), .B(
        Midori_rounds_SR_Result3[28]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[28]) );
  XNOR2_X1 Midori_rounds_U507 ( .A(Midori_rounds_SR_Result3[0]), .B(
        Midori_rounds_n1595), .ZN(Midori_rounds_n1445) );
  AOI22_X1 Midori_rounds_U506 ( .A1(Midori_rounds_n1274), .A2(Key3[28]), .B1(
        Key3[92]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1595) );
  MUX2_X1 Midori_rounds_U505 ( .A(Midori_rounds_n1444), .B(
        Midori_rounds_SR_Result3[27]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input3[27]) );
  XNOR2_X1 Midori_rounds_U504 ( .A(Midori_rounds_SR_Result3[31]), .B(
        Midori_rounds_n1598), .ZN(Midori_rounds_n1444) );
  AOI22_X1 Midori_rounds_U503 ( .A1(Midori_rounds_n1274), .A2(Key3[27]), .B1(
        Key3[91]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1598) );
  MUX2_X1 Midori_rounds_U502 ( .A(Midori_rounds_n1443), .B(
        Midori_rounds_SR_Result3[26]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input3[26]) );
  XNOR2_X1 Midori_rounds_U501 ( .A(Midori_rounds_SR_Result3[30]), .B(
        Midori_rounds_n1601), .ZN(Midori_rounds_n1443) );
  AOI22_X1 Midori_rounds_U500 ( .A1(Midori_rounds_n1274), .A2(Key3[26]), .B1(
        Key3[90]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1601) );
  MUX2_X1 Midori_rounds_U499 ( .A(Midori_rounds_n1442), .B(
        Midori_rounds_SR_Result3[25]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[25]) );
  XNOR2_X1 Midori_rounds_U498 ( .A(Midori_rounds_SR_Result3[29]), .B(
        Midori_rounds_n1604), .ZN(Midori_rounds_n1442) );
  AOI22_X1 Midori_rounds_U497 ( .A1(Midori_rounds_n1274), .A2(Key3[25]), .B1(
        Key3[89]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1604) );
  MUX2_X1 Midori_rounds_U496 ( .A(Midori_rounds_n1441), .B(
        Midori_rounds_SR_Result3[24]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input3[24]) );
  XNOR2_X1 Midori_rounds_U495 ( .A(Midori_rounds_SR_Result3[28]), .B(
        Midori_rounds_n1607), .ZN(Midori_rounds_n1441) );
  AOI22_X1 Midori_rounds_U494 ( .A1(Midori_rounds_n1274), .A2(Key3[24]), .B1(
        Key3[88]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1607) );
  MUX2_X1 Midori_rounds_U493 ( .A(Midori_rounds_n1440), .B(
        Midori_rounds_SR_Result3[23]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[23]) );
  XNOR2_X1 Midori_rounds_U492 ( .A(Midori_rounds_SR_Result3[59]), .B(
        Midori_rounds_n1610), .ZN(Midori_rounds_n1440) );
  AOI22_X1 Midori_rounds_U491 ( .A1(Midori_rounds_n1274), .A2(Key3[23]), .B1(
        Key3[87]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1610) );
  MUX2_X1 Midori_rounds_U490 ( .A(Midori_rounds_n1439), .B(
        Midori_rounds_SR_Result3[22]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[22]) );
  XNOR2_X1 Midori_rounds_U489 ( .A(Midori_rounds_SR_Result3[58]), .B(
        Midori_rounds_n1613), .ZN(Midori_rounds_n1439) );
  AOI22_X1 Midori_rounds_U488 ( .A1(Midori_rounds_n1274), .A2(Key3[22]), .B1(
        Key3[86]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1613) );
  MUX2_X1 Midori_rounds_U487 ( .A(Midori_rounds_n1438), .B(
        Midori_rounds_SR_Result3[21]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[21]) );
  XNOR2_X1 Midori_rounds_U486 ( .A(Midori_rounds_SR_Result3[57]), .B(
        Midori_rounds_n1616), .ZN(Midori_rounds_n1438) );
  AOI22_X1 Midori_rounds_U485 ( .A1(Midori_rounds_n1273), .A2(Key3[21]), .B1(
        Key3[85]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1616) );
  MUX2_X1 Midori_rounds_U484 ( .A(Midori_rounds_n1437), .B(
        Midori_rounds_SR_Result3[20]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[20]) );
  XNOR2_X1 Midori_rounds_U483 ( .A(Midori_rounds_SR_Result3[56]), .B(
        Midori_rounds_n1619), .ZN(Midori_rounds_n1437) );
  AOI22_X1 Midori_rounds_U482 ( .A1(Midori_rounds_n1273), .A2(Key3[20]), .B1(
        Key3[84]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1619) );
  MUX2_X1 Midori_rounds_U481 ( .A(Midori_rounds_n1436), .B(
        Midori_rounds_SR_Result3[1]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[1]) );
  XNOR2_X1 Midori_rounds_U480 ( .A(Midori_rounds_SR_Result3[49]), .B(
        Midori_rounds_n1676), .ZN(Midori_rounds_n1436) );
  AOI22_X1 Midori_rounds_U479 ( .A1(Midori_rounds_n1273), .A2(Key3[1]), .B1(
        Key3[65]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1676) );
  MUX2_X1 Midori_rounds_U478 ( .A(Midori_rounds_n1435), .B(
        Midori_rounds_SR_Result3[19]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[19]) );
  XNOR2_X1 Midori_rounds_U477 ( .A(Midori_rounds_SR_Result3[39]), .B(
        Midori_rounds_n1622), .ZN(Midori_rounds_n1435) );
  AOI22_X1 Midori_rounds_U476 ( .A1(Midori_rounds_n1273), .A2(Key3[19]), .B1(
        Key3[83]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1622) );
  MUX2_X1 Midori_rounds_U475 ( .A(Midori_rounds_n1434), .B(
        Midori_rounds_SR_Result3[18]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[18]) );
  XNOR2_X1 Midori_rounds_U474 ( .A(Midori_rounds_SR_Result3[38]), .B(
        Midori_rounds_n1625), .ZN(Midori_rounds_n1434) );
  AOI22_X1 Midori_rounds_U473 ( .A1(Midori_rounds_n1273), .A2(Key3[18]), .B1(
        Key3[82]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1625) );
  MUX2_X1 Midori_rounds_U472 ( .A(Midori_rounds_n1433), .B(
        Midori_rounds_SR_Result3[17]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[17]) );
  XNOR2_X1 Midori_rounds_U471 ( .A(Midori_rounds_SR_Result3[37]), .B(
        Midori_rounds_n1628), .ZN(Midori_rounds_n1433) );
  AOI22_X1 Midori_rounds_U470 ( .A1(Midori_rounds_n1273), .A2(Key3[17]), .B1(
        Key3[81]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1628) );
  MUX2_X1 Midori_rounds_U469 ( .A(Midori_rounds_n1432), .B(
        Midori_rounds_SR_Result3[16]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[16]) );
  XNOR2_X1 Midori_rounds_U468 ( .A(Midori_rounds_SR_Result3[36]), .B(
        Midori_rounds_n1631), .ZN(Midori_rounds_n1432) );
  AOI22_X1 Midori_rounds_U467 ( .A1(Midori_rounds_n1273), .A2(Key3[16]), .B1(
        Key3[80]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1631) );
  MUX2_X1 Midori_rounds_U466 ( .A(Midori_rounds_n1431), .B(
        Midori_rounds_SR_Result3[15]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[15]) );
  XNOR2_X1 Midori_rounds_U465 ( .A(Midori_rounds_SR_Result3[23]), .B(
        Midori_rounds_n1634), .ZN(Midori_rounds_n1431) );
  AOI22_X1 Midori_rounds_U464 ( .A1(Midori_rounds_n1273), .A2(Key3[15]), .B1(
        Key3[79]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1634) );
  MUX2_X1 Midori_rounds_U463 ( .A(Midori_rounds_n1430), .B(
        Midori_rounds_SR_Result3[14]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[14]) );
  XNOR2_X1 Midori_rounds_U462 ( .A(Midori_rounds_SR_Result3[22]), .B(
        Midori_rounds_n1637), .ZN(Midori_rounds_n1430) );
  AOI22_X1 Midori_rounds_U461 ( .A1(Midori_rounds_n1273), .A2(Key3[14]), .B1(
        Key3[78]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1637) );
  MUX2_X1 Midori_rounds_U460 ( .A(Midori_rounds_n1429), .B(
        Midori_rounds_SR_Result3[13]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input3[13]) );
  XNOR2_X1 Midori_rounds_U459 ( .A(Midori_rounds_SR_Result3[21]), .B(
        Midori_rounds_n1640), .ZN(Midori_rounds_n1429) );
  AOI22_X1 Midori_rounds_U458 ( .A1(Midori_rounds_n1273), .A2(Key3[13]), .B1(
        Key3[77]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1640) );
  MUX2_X1 Midori_rounds_U457 ( .A(Midori_rounds_n1428), .B(
        Midori_rounds_SR_Result3[12]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input3[12]) );
  XNOR2_X1 Midori_rounds_U456 ( .A(Midori_rounds_SR_Result3[20]), .B(
        Midori_rounds_n1643), .ZN(Midori_rounds_n1428) );
  AOI22_X1 Midori_rounds_U455 ( .A1(Midori_rounds_n1273), .A2(Key3[12]), .B1(
        Key3[76]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1643) );
  MUX2_X1 Midori_rounds_U454 ( .A(Midori_rounds_n1427), .B(
        Midori_rounds_SR_Result3[11]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[11]) );
  XNOR2_X1 Midori_rounds_U453 ( .A(Midori_rounds_SR_Result3[11]), .B(
        Midori_rounds_n1646), .ZN(Midori_rounds_n1427) );
  AOI22_X1 Midori_rounds_U452 ( .A1(Midori_rounds_n1273), .A2(Key3[11]), .B1(
        Key3[75]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1646) );
  MUX2_X1 Midori_rounds_U451 ( .A(Midori_rounds_n1426), .B(
        Midori_rounds_SR_Result3[10]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input3[10]) );
  XNOR2_X1 Midori_rounds_U450 ( .A(Midori_rounds_SR_Result3[10]), .B(
        Midori_rounds_n1649), .ZN(Midori_rounds_n1426) );
  AOI22_X1 Midori_rounds_U449 ( .A1(Midori_rounds_n1273), .A2(Key3[10]), .B1(
        Key3[74]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1649) );
  MUX2_X1 Midori_rounds_U448 ( .A(Midori_rounds_n1425), .B(
        Midori_rounds_SR_Result3[0]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input3[0]) );
  XNOR2_X1 Midori_rounds_U447 ( .A(Midori_rounds_SR_Result3[48]), .B(
        Midori_rounds_n1679), .ZN(Midori_rounds_n1425) );
  AOI22_X1 Midori_rounds_U446 ( .A1(Midori_rounds_n1272), .A2(Key3[0]), .B1(
        Key3[64]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1679) );
  MUX2_X1 Midori_rounds_U445 ( .A(Midori_rounds_n1424), .B(
        Midori_rounds_SR_Result2[9]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input2[9]) );
  XNOR2_X1 Midori_rounds_U444 ( .A(Midori_rounds_SR_Result2[9]), .B(
        Midori_rounds_n1844), .ZN(Midori_rounds_n1424) );
  AOI22_X1 Midori_rounds_U443 ( .A1(Midori_rounds_n1272), .A2(Key2[9]), .B1(
        Key2[73]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1844) );
  MUX2_X1 Midori_rounds_U442 ( .A(Midori_rounds_n1423), .B(
        Midori_rounds_SR_Result2[8]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input2[8]) );
  XNOR2_X1 Midori_rounds_U441 ( .A(Midori_rounds_SR_Result2[8]), .B(
        Midori_rounds_n1847), .ZN(Midori_rounds_n1423) );
  AOI22_X1 Midori_rounds_U440 ( .A1(Midori_rounds_n1272), .A2(Key2[8]), .B1(
        Key2[72]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1847) );
  MUX2_X1 Midori_rounds_U439 ( .A(Midori_rounds_n1422), .B(
        Midori_rounds_SR_Result2[7]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input2[7]) );
  XNOR2_X1 Midori_rounds_U438 ( .A(Midori_rounds_SR_Result2[47]), .B(
        Midori_rounds_n1850), .ZN(Midori_rounds_n1422) );
  AOI22_X1 Midori_rounds_U437 ( .A1(Midori_rounds_n1272), .A2(Key2[7]), .B1(
        Key2[71]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1850) );
  MUX2_X1 Midori_rounds_U436 ( .A(Midori_rounds_n1421), .B(
        Midori_rounds_SR_Result2[6]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input2[6]) );
  XNOR2_X1 Midori_rounds_U435 ( .A(Midori_rounds_SR_Result2[46]), .B(
        Midori_rounds_n1853), .ZN(Midori_rounds_n1421) );
  AOI22_X1 Midori_rounds_U434 ( .A1(Midori_rounds_n1272), .A2(Key2[6]), .B1(
        Key2[70]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1853) );
  MUX2_X1 Midori_rounds_U433 ( .A(Midori_rounds_n1420), .B(
        Midori_rounds_SR_Result2[63]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input2[63]) );
  XNOR2_X1 Midori_rounds_U432 ( .A(Midori_rounds_SR_Result2[63]), .B(
        Midori_rounds_n1682), .ZN(Midori_rounds_n1420) );
  AOI22_X1 Midori_rounds_U431 ( .A1(Midori_rounds_n1272), .A2(Key2[63]), .B1(
        Key2[127]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1682) );
  MUX2_X1 Midori_rounds_U430 ( .A(Midori_rounds_n1419), .B(
        Midori_rounds_SR_Result2[62]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input2[62]) );
  XNOR2_X1 Midori_rounds_U429 ( .A(Midori_rounds_SR_Result2[62]), .B(
        Midori_rounds_n1685), .ZN(Midori_rounds_n1419) );
  AOI22_X1 Midori_rounds_U428 ( .A1(Midori_rounds_n1272), .A2(Key2[62]), .B1(
        Key2[126]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1685) );
  MUX2_X1 Midori_rounds_U427 ( .A(Midori_rounds_n1418), .B(
        Midori_rounds_SR_Result2[61]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input2[61]) );
  XNOR2_X1 Midori_rounds_U426 ( .A(Midori_rounds_SR_Result2[61]), .B(
        Midori_rounds_n1688), .ZN(Midori_rounds_n1418) );
  AOI22_X1 Midori_rounds_U425 ( .A1(Midori_rounds_n1272), .A2(Key2[61]), .B1(
        Key2[125]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1688) );
  MUX2_X1 Midori_rounds_U424 ( .A(Midori_rounds_n1417), .B(
        Midori_rounds_SR_Result2[60]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input2[60]) );
  XNOR2_X1 Midori_rounds_U423 ( .A(Midori_rounds_SR_Result2[60]), .B(
        Midori_rounds_n1691), .ZN(Midori_rounds_n1417) );
  AOI22_X1 Midori_rounds_U422 ( .A1(Midori_rounds_n1272), .A2(Key2[60]), .B1(
        Key2[124]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1691) );
  MUX2_X1 Midori_rounds_U421 ( .A(Midori_rounds_n1416), .B(
        Midori_rounds_SR_Result2[5]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input2[5]) );
  XNOR2_X1 Midori_rounds_U420 ( .A(Midori_rounds_SR_Result2[45]), .B(
        Midori_rounds_n1856), .ZN(Midori_rounds_n1416) );
  AOI22_X1 Midori_rounds_U419 ( .A1(Midori_rounds_n1272), .A2(Key2[5]), .B1(
        Key2[69]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1856) );
  MUX2_X1 Midori_rounds_U418 ( .A(Midori_rounds_n1415), .B(
        Midori_rounds_SR_Result2[59]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input2[59]) );
  XNOR2_X1 Midori_rounds_U417 ( .A(Midori_rounds_SR_Result2[35]), .B(
        Midori_rounds_n1694), .ZN(Midori_rounds_n1415) );
  AOI22_X1 Midori_rounds_U416 ( .A1(Midori_rounds_n1272), .A2(Key2[59]), .B1(
        Key2[123]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1694) );
  MUX2_X1 Midori_rounds_U415 ( .A(Midori_rounds_n1414), .B(
        Midori_rounds_SR_Result2[58]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input2[58]) );
  XNOR2_X1 Midori_rounds_U414 ( .A(Midori_rounds_SR_Result2[34]), .B(
        Midori_rounds_n1697), .ZN(Midori_rounds_n1414) );
  AOI22_X1 Midori_rounds_U413 ( .A1(Midori_rounds_n1272), .A2(Key2[58]), .B1(
        Key2[122]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1697) );
  MUX2_X1 Midori_rounds_U412 ( .A(Midori_rounds_n1413), .B(
        Midori_rounds_SR_Result2[57]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input2[57]) );
  XNOR2_X1 Midori_rounds_U411 ( .A(Midori_rounds_SR_Result2[33]), .B(
        Midori_rounds_n1700), .ZN(Midori_rounds_n1413) );
  AOI22_X1 Midori_rounds_U410 ( .A1(Midori_rounds_n1272), .A2(Key2[57]), .B1(
        Key2[121]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1700) );
  MUX2_X1 Midori_rounds_U409 ( .A(Midori_rounds_n1412), .B(
        Midori_rounds_SR_Result2[56]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input2[56]) );
  XNOR2_X1 Midori_rounds_U408 ( .A(Midori_rounds_SR_Result2[32]), .B(
        Midori_rounds_n1703), .ZN(Midori_rounds_n1412) );
  AOI22_X1 Midori_rounds_U407 ( .A1(Midori_rounds_n1271), .A2(Key2[56]), .B1(
        Key2[120]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1703) );
  MUX2_X1 Midori_rounds_U406 ( .A(Midori_rounds_n1411), .B(
        Midori_rounds_SR_Result2[55]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input2[55]) );
  XNOR2_X1 Midori_rounds_U405 ( .A(Midori_rounds_SR_Result2[7]), .B(
        Midori_rounds_n1706), .ZN(Midori_rounds_n1411) );
  AOI22_X1 Midori_rounds_U404 ( .A1(Midori_rounds_n1271), .A2(Key2[55]), .B1(
        Key2[119]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1706) );
  MUX2_X1 Midori_rounds_U403 ( .A(Midori_rounds_n1410), .B(
        Midori_rounds_SR_Result2[54]), .S(Midori_rounds_n1245), .Z(
        Midori_rounds_mul_input2[54]) );
  XNOR2_X1 Midori_rounds_U402 ( .A(Midori_rounds_SR_Result2[6]), .B(
        Midori_rounds_n1709), .ZN(Midori_rounds_n1410) );
  AOI22_X1 Midori_rounds_U401 ( .A1(Midori_rounds_n1271), .A2(Key2[54]), .B1(
        Key2[118]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1709) );
  MUX2_X1 Midori_rounds_U400 ( .A(Midori_rounds_n1409), .B(
        Midori_rounds_SR_Result2[53]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input2[53]) );
  XNOR2_X1 Midori_rounds_U399 ( .A(Midori_rounds_SR_Result2[5]), .B(
        Midori_rounds_n1712), .ZN(Midori_rounds_n1409) );
  AOI22_X1 Midori_rounds_U398 ( .A1(Midori_rounds_n1271), .A2(Key2[53]), .B1(
        Key2[117]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1712) );
  MUX2_X1 Midori_rounds_U397 ( .A(Midori_rounds_n1408), .B(
        Midori_rounds_SR_Result2[52]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input2[52]) );
  XNOR2_X1 Midori_rounds_U396 ( .A(Midori_rounds_SR_Result2[4]), .B(
        Midori_rounds_n1715), .ZN(Midori_rounds_n1408) );
  AOI22_X1 Midori_rounds_U395 ( .A1(Midori_rounds_n1271), .A2(Key2[52]), .B1(
        Key2[116]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1715) );
  MUX2_X1 Midori_rounds_U394 ( .A(Midori_rounds_n1407), .B(
        Midori_rounds_SR_Result2[51]), .S(Midori_rounds_n1490), .Z(
        Midori_rounds_mul_input2[51]) );
  XNOR2_X1 Midori_rounds_U393 ( .A(Midori_rounds_SR_Result2[27]), .B(
        Midori_rounds_n1718), .ZN(Midori_rounds_n1407) );
  AOI22_X1 Midori_rounds_U392 ( .A1(Midori_rounds_n1271), .A2(Key2[51]), .B1(
        Key2[115]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1718) );
  MUX2_X1 Midori_rounds_U391 ( .A(Midori_rounds_n1406), .B(
        Midori_rounds_SR_Result2[50]), .S(Midori_rounds_n1246), .Z(
        Midori_rounds_mul_input2[50]) );
  XNOR2_X1 Midori_rounds_U390 ( .A(Midori_rounds_SR_Result2[26]), .B(
        Midori_rounds_n1721), .ZN(Midori_rounds_n1406) );
  AOI22_X1 Midori_rounds_U389 ( .A1(Midori_rounds_n1271), .A2(Key2[50]), .B1(
        Key2[114]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1721) );
  MUX2_X1 Midori_rounds_U388 ( .A(Midori_rounds_n1405), .B(
        Midori_rounds_SR_Result2[4]), .S(Midori_rounds_n1250), .Z(
        Midori_rounds_mul_input2[4]) );
  XNOR2_X1 Midori_rounds_U387 ( .A(Midori_rounds_SR_Result2[44]), .B(
        Midori_rounds_n1859), .ZN(Midori_rounds_n1405) );
  AOI22_X1 Midori_rounds_U386 ( .A1(Midori_rounds_n1271), .A2(Key2[4]), .B1(
        Key2[68]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1859) );
  MUX2_X1 Midori_rounds_U385 ( .A(Midori_rounds_n1404), .B(
        Midori_rounds_SR_Result2[49]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[49]) );
  XNOR2_X1 Midori_rounds_U384 ( .A(Midori_rounds_SR_Result2[25]), .B(
        Midori_rounds_n1724), .ZN(Midori_rounds_n1404) );
  AOI22_X1 Midori_rounds_U383 ( .A1(Midori_rounds_n1271), .A2(Key2[49]), .B1(
        Key2[113]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1724) );
  MUX2_X1 Midori_rounds_U382 ( .A(Midori_rounds_n1403), .B(
        Midori_rounds_SR_Result2[48]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[48]) );
  XNOR2_X1 Midori_rounds_U381 ( .A(Midori_rounds_SR_Result2[24]), .B(
        Midori_rounds_n1727), .ZN(Midori_rounds_n1403) );
  AOI22_X1 Midori_rounds_U380 ( .A1(Midori_rounds_n1271), .A2(Key2[48]), .B1(
        Key2[112]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1727) );
  MUX2_X1 Midori_rounds_U379 ( .A(Midori_rounds_n1402), .B(
        Midori_rounds_SR_Result2[47]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[47]) );
  XNOR2_X1 Midori_rounds_U378 ( .A(Midori_rounds_SR_Result2[43]), .B(
        Midori_rounds_n1730), .ZN(Midori_rounds_n1402) );
  AOI22_X1 Midori_rounds_U377 ( .A1(Midori_rounds_n1271), .A2(Key2[47]), .B1(
        Key2[111]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1730) );
  MUX2_X1 Midori_rounds_U376 ( .A(Midori_rounds_n1401), .B(
        Midori_rounds_SR_Result2[46]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[46]) );
  XNOR2_X1 Midori_rounds_U375 ( .A(Midori_rounds_SR_Result2[42]), .B(
        Midori_rounds_n1733), .ZN(Midori_rounds_n1401) );
  AOI22_X1 Midori_rounds_U374 ( .A1(Midori_rounds_n1271), .A2(Key2[46]), .B1(
        Key2[110]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1733) );
  MUX2_X1 Midori_rounds_U373 ( .A(Midori_rounds_n1400), .B(
        Midori_rounds_SR_Result2[45]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[45]) );
  XNOR2_X1 Midori_rounds_U372 ( .A(Midori_rounds_SR_Result2[41]), .B(
        Midori_rounds_n1736), .ZN(Midori_rounds_n1400) );
  AOI22_X1 Midori_rounds_U371 ( .A1(Midori_rounds_n1271), .A2(Key2[45]), .B1(
        Key2[109]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1736) );
  MUX2_X1 Midori_rounds_U370 ( .A(Midori_rounds_n1399), .B(
        Midori_rounds_SR_Result2[44]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[44]) );
  XNOR2_X1 Midori_rounds_U369 ( .A(Midori_rounds_SR_Result2[40]), .B(
        Midori_rounds_n1739), .ZN(Midori_rounds_n1399) );
  AOI22_X1 Midori_rounds_U368 ( .A1(Midori_rounds_n1270), .A2(Key2[44]), .B1(
        Key2[108]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1739) );
  MUX2_X1 Midori_rounds_U367 ( .A(Midori_rounds_n1398), .B(
        Midori_rounds_SR_Result2[43]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[43]) );
  XNOR2_X1 Midori_rounds_U366 ( .A(Midori_rounds_SR_Result2[55]), .B(
        Midori_rounds_n1742), .ZN(Midori_rounds_n1398) );
  AOI22_X1 Midori_rounds_U365 ( .A1(Midori_rounds_n1270), .A2(Key2[43]), .B1(
        Key2[107]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1742) );
  MUX2_X1 Midori_rounds_U364 ( .A(Midori_rounds_n1397), .B(
        Midori_rounds_SR_Result2[42]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[42]) );
  XNOR2_X1 Midori_rounds_U363 ( .A(Midori_rounds_SR_Result2[54]), .B(
        Midori_rounds_n1745), .ZN(Midori_rounds_n1397) );
  AOI22_X1 Midori_rounds_U362 ( .A1(Midori_rounds_n1270), .A2(Key2[42]), .B1(
        Key2[106]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1745) );
  MUX2_X1 Midori_rounds_U361 ( .A(Midori_rounds_n1396), .B(
        Midori_rounds_SR_Result2[41]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[41]) );
  XNOR2_X1 Midori_rounds_U360 ( .A(Midori_rounds_SR_Result2[53]), .B(
        Midori_rounds_n1748), .ZN(Midori_rounds_n1396) );
  AOI22_X1 Midori_rounds_U359 ( .A1(Midori_rounds_n1270), .A2(Key2[41]), .B1(
        Key2[105]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1748) );
  MUX2_X1 Midori_rounds_U358 ( .A(Midori_rounds_n1395), .B(
        Midori_rounds_SR_Result2[40]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[40]) );
  XNOR2_X1 Midori_rounds_U357 ( .A(Midori_rounds_SR_Result2[52]), .B(
        Midori_rounds_n1751), .ZN(Midori_rounds_n1395) );
  AOI22_X1 Midori_rounds_U356 ( .A1(Midori_rounds_n1270), .A2(Key2[40]), .B1(
        Key2[104]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1751) );
  MUX2_X1 Midori_rounds_U355 ( .A(Midori_rounds_n1394), .B(
        Midori_rounds_SR_Result2[3]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[3]) );
  XNOR2_X1 Midori_rounds_U354 ( .A(Midori_rounds_SR_Result2[51]), .B(
        Midori_rounds_n1862), .ZN(Midori_rounds_n1394) );
  AOI22_X1 Midori_rounds_U353 ( .A1(Midori_rounds_n1270), .A2(Key2[3]), .B1(
        Key2[67]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1862) );
  MUX2_X1 Midori_rounds_U352 ( .A(Midori_rounds_n1393), .B(
        Midori_rounds_SR_Result2[39]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[39]) );
  XNOR2_X1 Midori_rounds_U351 ( .A(Midori_rounds_SR_Result2[19]), .B(
        Midori_rounds_n1754), .ZN(Midori_rounds_n1393) );
  AOI22_X1 Midori_rounds_U350 ( .A1(Midori_rounds_n1270), .A2(Key2[39]), .B1(
        Key2[103]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1754) );
  MUX2_X1 Midori_rounds_U349 ( .A(Midori_rounds_n1392), .B(
        Midori_rounds_SR_Result2[38]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[38]) );
  XNOR2_X1 Midori_rounds_U348 ( .A(Midori_rounds_SR_Result2[18]), .B(
        Midori_rounds_n1757), .ZN(Midori_rounds_n1392) );
  AOI22_X1 Midori_rounds_U347 ( .A1(Midori_rounds_n1270), .A2(Key2[38]), .B1(
        Key2[102]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1757) );
  MUX2_X1 Midori_rounds_U346 ( .A(Midori_rounds_n1391), .B(
        Midori_rounds_SR_Result2[37]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[37]) );
  XNOR2_X1 Midori_rounds_U345 ( .A(Midori_rounds_SR_Result2[17]), .B(
        Midori_rounds_n1760), .ZN(Midori_rounds_n1391) );
  AOI22_X1 Midori_rounds_U344 ( .A1(Midori_rounds_n1270), .A2(Key2[37]), .B1(
        Key2[101]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1760) );
  MUX2_X1 Midori_rounds_U343 ( .A(Midori_rounds_n1390), .B(
        Midori_rounds_SR_Result2[36]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[36]) );
  XNOR2_X1 Midori_rounds_U342 ( .A(Midori_rounds_SR_Result2[16]), .B(
        Midori_rounds_n1763), .ZN(Midori_rounds_n1390) );
  AOI22_X1 Midori_rounds_U341 ( .A1(Midori_rounds_n1270), .A2(Key2[36]), .B1(
        Key2[100]), .B2(Midori_rounds_n1280), .ZN(Midori_rounds_n1763) );
  MUX2_X1 Midori_rounds_U340 ( .A(Midori_rounds_n1389), .B(
        Midori_rounds_SR_Result2[35]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[35]) );
  XNOR2_X1 Midori_rounds_U339 ( .A(Midori_rounds_SR_Result2[15]), .B(
        Midori_rounds_n1766), .ZN(Midori_rounds_n1389) );
  AOI22_X1 Midori_rounds_U338 ( .A1(Midori_rounds_n1270), .A2(Key2[35]), .B1(
        Key2[99]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1766) );
  MUX2_X1 Midori_rounds_U337 ( .A(Midori_rounds_n1388), .B(
        Midori_rounds_SR_Result2[34]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[34]) );
  XNOR2_X1 Midori_rounds_U336 ( .A(Midori_rounds_SR_Result2[14]), .B(
        Midori_rounds_n1769), .ZN(Midori_rounds_n1388) );
  AOI22_X1 Midori_rounds_U335 ( .A1(Midori_rounds_n1270), .A2(Key2[34]), .B1(
        Key2[98]), .B2(Midori_rounds_n1275), .ZN(Midori_rounds_n1769) );
  MUX2_X1 Midori_rounds_U334 ( .A(Midori_rounds_n1387), .B(
        Midori_rounds_SR_Result2[33]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[33]) );
  XNOR2_X1 Midori_rounds_U333 ( .A(Midori_rounds_SR_Result2[13]), .B(
        Midori_rounds_n1772), .ZN(Midori_rounds_n1387) );
  AOI22_X1 Midori_rounds_U332 ( .A1(Midori_rounds_n1270), .A2(Key2[33]), .B1(
        Key2[97]), .B2(Midori_rounds_n1275), .ZN(Midori_rounds_n1772) );
  MUX2_X1 Midori_rounds_U331 ( .A(Midori_rounds_n1386), .B(
        Midori_rounds_SR_Result2[32]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[32]) );
  XNOR2_X1 Midori_rounds_U330 ( .A(Midori_rounds_SR_Result2[12]), .B(
        Midori_rounds_n1775), .ZN(Midori_rounds_n1386) );
  AOI22_X1 Midori_rounds_U329 ( .A1(Midori_rounds_n1270), .A2(Key2[32]), .B1(
        Key2[96]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1775) );
  MUX2_X1 Midori_rounds_U328 ( .A(Midori_rounds_n1385), .B(
        Midori_rounds_SR_Result2[31]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[31]) );
  XNOR2_X1 Midori_rounds_U327 ( .A(Midori_rounds_SR_Result2[3]), .B(
        Midori_rounds_n1778), .ZN(Midori_rounds_n1385) );
  AOI22_X1 Midori_rounds_U326 ( .A1(Midori_rounds_n1273), .A2(Key2[31]), .B1(
        Key2[95]), .B2(Midori_rounds_n1275), .ZN(Midori_rounds_n1778) );
  MUX2_X1 Midori_rounds_U325 ( .A(Midori_rounds_n1384), .B(
        Midori_rounds_SR_Result2[30]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[30]) );
  XNOR2_X1 Midori_rounds_U324 ( .A(Midori_rounds_SR_Result2[2]), .B(
        Midori_rounds_n1781), .ZN(Midori_rounds_n1384) );
  AOI22_X1 Midori_rounds_U323 ( .A1(Midori_rounds_n1269), .A2(Key2[30]), .B1(
        Key2[94]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1781) );
  MUX2_X1 Midori_rounds_U322 ( .A(Midori_rounds_n1383), .B(
        Midori_rounds_SR_Result2[2]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[2]) );
  XNOR2_X1 Midori_rounds_U321 ( .A(Midori_rounds_SR_Result2[50]), .B(
        Midori_rounds_n1865), .ZN(Midori_rounds_n1383) );
  AOI22_X1 Midori_rounds_U320 ( .A1(Midori_rounds_n1272), .A2(Key2[2]), .B1(
        Key2[66]), .B2(Midori_rounds_n1275), .ZN(Midori_rounds_n1865) );
  MUX2_X1 Midori_rounds_U319 ( .A(Midori_rounds_n1382), .B(
        Midori_rounds_SR_Result2[29]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[29]) );
  XNOR2_X1 Midori_rounds_U318 ( .A(Midori_rounds_SR_Result2[1]), .B(
        Midori_rounds_n1784), .ZN(Midori_rounds_n1382) );
  AOI22_X1 Midori_rounds_U317 ( .A1(Midori_rounds_n1273), .A2(Key2[29]), .B1(
        Key2[93]), .B2(Midori_rounds_n1275), .ZN(Midori_rounds_n1784) );
  MUX2_X1 Midori_rounds_U316 ( .A(Midori_rounds_n1381), .B(
        Midori_rounds_SR_Result2[28]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[28]) );
  XNOR2_X1 Midori_rounds_U315 ( .A(Midori_rounds_SR_Result2[0]), .B(
        Midori_rounds_n1787), .ZN(Midori_rounds_n1381) );
  AOI22_X1 Midori_rounds_U314 ( .A1(Midori_rounds_n1272), .A2(Key2[28]), .B1(
        Key2[92]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1787) );
  MUX2_X1 Midori_rounds_U313 ( .A(Midori_rounds_n1380), .B(
        Midori_rounds_SR_Result2[27]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[27]) );
  XNOR2_X1 Midori_rounds_U312 ( .A(Midori_rounds_SR_Result2[31]), .B(
        Midori_rounds_n1790), .ZN(Midori_rounds_n1380) );
  AOI22_X1 Midori_rounds_U311 ( .A1(Midori_rounds_n1271), .A2(Key2[27]), .B1(
        Key2[91]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1790) );
  MUX2_X1 Midori_rounds_U310 ( .A(Midori_rounds_n1379), .B(
        Midori_rounds_SR_Result2[26]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[26]) );
  XNOR2_X1 Midori_rounds_U309 ( .A(Midori_rounds_SR_Result2[30]), .B(
        Midori_rounds_n1793), .ZN(Midori_rounds_n1379) );
  AOI22_X1 Midori_rounds_U308 ( .A1(Midori_rounds_n1273), .A2(Key2[26]), .B1(
        Key2[90]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1793) );
  MUX2_X1 Midori_rounds_U307 ( .A(Midori_rounds_n1378), .B(
        Midori_rounds_SR_Result2[25]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[25]) );
  XNOR2_X1 Midori_rounds_U306 ( .A(Midori_rounds_SR_Result2[29]), .B(
        Midori_rounds_n1796), .ZN(Midori_rounds_n1378) );
  AOI22_X1 Midori_rounds_U305 ( .A1(Midori_rounds_n1270), .A2(Key2[25]), .B1(
        Key2[89]), .B2(Midori_rounds_n1275), .ZN(Midori_rounds_n1796) );
  MUX2_X1 Midori_rounds_U304 ( .A(Midori_rounds_n1377), .B(
        Midori_rounds_SR_Result2[24]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[24]) );
  XNOR2_X1 Midori_rounds_U303 ( .A(Midori_rounds_SR_Result2[28]), .B(
        Midori_rounds_n1799), .ZN(Midori_rounds_n1377) );
  AOI22_X1 Midori_rounds_U302 ( .A1(Midori_rounds_n1271), .A2(Key2[24]), .B1(
        Key2[88]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1799) );
  MUX2_X1 Midori_rounds_U301 ( .A(Midori_rounds_n1376), .B(
        Midori_rounds_SR_Result2[23]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[23]) );
  XNOR2_X1 Midori_rounds_U300 ( .A(Midori_rounds_SR_Result2[59]), .B(
        Midori_rounds_n1802), .ZN(Midori_rounds_n1376) );
  AOI22_X1 Midori_rounds_U299 ( .A1(Midori_rounds_n1272), .A2(Key2[23]), .B1(
        Key2[87]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1802) );
  MUX2_X1 Midori_rounds_U298 ( .A(Midori_rounds_n1375), .B(
        Midori_rounds_SR_Result2[22]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[22]) );
  XNOR2_X1 Midori_rounds_U297 ( .A(Midori_rounds_SR_Result2[58]), .B(
        Midori_rounds_n1805), .ZN(Midori_rounds_n1375) );
  AOI22_X1 Midori_rounds_U296 ( .A1(Midori_rounds_n1274), .A2(Key2[22]), .B1(
        Key2[86]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1805) );
  MUX2_X1 Midori_rounds_U295 ( .A(Midori_rounds_n1374), .B(
        Midori_rounds_SR_Result2[21]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[21]) );
  XNOR2_X1 Midori_rounds_U294 ( .A(Midori_rounds_SR_Result2[57]), .B(
        Midori_rounds_n1808), .ZN(Midori_rounds_n1374) );
  AOI22_X1 Midori_rounds_U293 ( .A1(Midori_rounds_n1274), .A2(Key2[21]), .B1(
        Key2[85]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1808) );
  MUX2_X1 Midori_rounds_U292 ( .A(Midori_rounds_n1373), .B(
        Midori_rounds_SR_Result2[20]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[20]) );
  XNOR2_X1 Midori_rounds_U291 ( .A(Midori_rounds_SR_Result2[56]), .B(
        Midori_rounds_n1811), .ZN(Midori_rounds_n1373) );
  AOI22_X1 Midori_rounds_U290 ( .A1(Midori_rounds_n1268), .A2(Key2[20]), .B1(
        Key2[84]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1811) );
  MUX2_X1 Midori_rounds_U289 ( .A(Midori_rounds_n1372), .B(
        Midori_rounds_SR_Result2[1]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[1]) );
  XNOR2_X1 Midori_rounds_U288 ( .A(Midori_rounds_SR_Result2[49]), .B(
        Midori_rounds_n1868), .ZN(Midori_rounds_n1372) );
  AOI22_X1 Midori_rounds_U287 ( .A1(Midori_rounds_n1270), .A2(Key2[1]), .B1(
        Key2[65]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1868) );
  MUX2_X1 Midori_rounds_U286 ( .A(Midori_rounds_n1371), .B(
        Midori_rounds_SR_Result2[19]), .S(Midori_rounds_n1247), .Z(
        Midori_rounds_mul_input2[19]) );
  XNOR2_X1 Midori_rounds_U285 ( .A(Midori_rounds_SR_Result2[39]), .B(
        Midori_rounds_n1814), .ZN(Midori_rounds_n1371) );
  AOI22_X1 Midori_rounds_U284 ( .A1(Midori_rounds_n1274), .A2(Key2[19]), .B1(
        Key2[83]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1814) );
  MUX2_X1 Midori_rounds_U283 ( .A(Midori_rounds_n1370), .B(
        Midori_rounds_SR_Result2[18]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[18]) );
  XNOR2_X1 Midori_rounds_U282 ( .A(Midori_rounds_SR_Result2[38]), .B(
        Midori_rounds_n1817), .ZN(Midori_rounds_n1370) );
  AOI22_X1 Midori_rounds_U281 ( .A1(Midori_rounds_n1273), .A2(Key2[18]), .B1(
        Key2[82]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1817) );
  MUX2_X1 Midori_rounds_U280 ( .A(Midori_rounds_n1369), .B(
        Midori_rounds_SR_Result2[17]), .S(Midori_rounds_n1244), .Z(
        Midori_rounds_mul_input2[17]) );
  XNOR2_X1 Midori_rounds_U279 ( .A(Midori_rounds_SR_Result2[37]), .B(
        Midori_rounds_n1820), .ZN(Midori_rounds_n1369) );
  AOI22_X1 Midori_rounds_U278 ( .A1(Midori_rounds_n1271), .A2(Key2[17]), .B1(
        Key2[81]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1820) );
  MUX2_X1 Midori_rounds_U277 ( .A(Midori_rounds_n1368), .B(
        Midori_rounds_SR_Result2[16]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input2[16]) );
  XNOR2_X1 Midori_rounds_U276 ( .A(Midori_rounds_SR_Result2[36]), .B(
        Midori_rounds_n1823), .ZN(Midori_rounds_n1368) );
  AOI22_X1 Midori_rounds_U275 ( .A1(Midori_rounds_n1273), .A2(Key2[16]), .B1(
        Key2[80]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1823) );
  MUX2_X1 Midori_rounds_U274 ( .A(Midori_rounds_n1367), .B(
        Midori_rounds_SR_Result2[15]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input2[15]) );
  XNOR2_X1 Midori_rounds_U273 ( .A(Midori_rounds_SR_Result2[23]), .B(
        Midori_rounds_n1826), .ZN(Midori_rounds_n1367) );
  AOI22_X1 Midori_rounds_U272 ( .A1(Midori_rounds_n1269), .A2(Key2[15]), .B1(
        Key2[79]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1826) );
  MUX2_X1 Midori_rounds_U271 ( .A(Midori_rounds_n1366), .B(
        Midori_rounds_SR_Result2[14]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input2[14]) );
  XNOR2_X1 Midori_rounds_U270 ( .A(Midori_rounds_SR_Result2[22]), .B(
        Midori_rounds_n1829), .ZN(Midori_rounds_n1366) );
  AOI22_X1 Midori_rounds_U269 ( .A1(Midori_rounds_n1274), .A2(Key2[14]), .B1(
        Key2[78]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1829) );
  MUX2_X1 Midori_rounds_U268 ( .A(Midori_rounds_n1365), .B(
        Midori_rounds_SR_Result2[13]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input2[13]) );
  XNOR2_X1 Midori_rounds_U267 ( .A(Midori_rounds_SR_Result2[21]), .B(
        Midori_rounds_n1832), .ZN(Midori_rounds_n1365) );
  AOI22_X1 Midori_rounds_U266 ( .A1(Midori_rounds_n1271), .A2(Key2[13]), .B1(
        Key2[77]), .B2(Midori_rounds_n1275), .ZN(Midori_rounds_n1832) );
  MUX2_X1 Midori_rounds_U265 ( .A(Midori_rounds_n1364), .B(
        Midori_rounds_SR_Result2[12]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input2[12]) );
  XNOR2_X1 Midori_rounds_U264 ( .A(Midori_rounds_SR_Result2[20]), .B(
        Midori_rounds_n1835), .ZN(Midori_rounds_n1364) );
  AOI22_X1 Midori_rounds_U263 ( .A1(Midori_rounds_n1270), .A2(Key2[12]), .B1(
        Key2[76]), .B2(Midori_rounds_n1275), .ZN(Midori_rounds_n1835) );
  MUX2_X1 Midori_rounds_U262 ( .A(Midori_rounds_n1363), .B(
        Midori_rounds_SR_Result2[11]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input2[11]) );
  XNOR2_X1 Midori_rounds_U261 ( .A(Midori_rounds_SR_Result2[11]), .B(
        Midori_rounds_n1838), .ZN(Midori_rounds_n1363) );
  AOI22_X1 Midori_rounds_U260 ( .A1(Midori_rounds_n1270), .A2(Key2[11]), .B1(
        Key2[75]), .B2(Midori_rounds_n1275), .ZN(Midori_rounds_n1838) );
  MUX2_X1 Midori_rounds_U259 ( .A(Midori_rounds_n1362), .B(
        Midori_rounds_SR_Result2[10]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input2[10]) );
  XNOR2_X1 Midori_rounds_U258 ( .A(Midori_rounds_SR_Result2[10]), .B(
        Midori_rounds_n1841), .ZN(Midori_rounds_n1362) );
  AOI22_X1 Midori_rounds_U257 ( .A1(Midori_rounds_n1271), .A2(Key2[10]), .B1(
        Key2[74]), .B2(Midori_rounds_n1275), .ZN(Midori_rounds_n1841) );
  MUX2_X1 Midori_rounds_U256 ( .A(Midori_rounds_n1361), .B(
        Midori_rounds_SR_Result2[0]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input2[0]) );
  XNOR2_X1 Midori_rounds_U255 ( .A(Midori_rounds_SR_Result2[48]), .B(
        Midori_rounds_n1871), .ZN(Midori_rounds_n1361) );
  AOI22_X1 Midori_rounds_U254 ( .A1(Midori_rounds_n1274), .A2(Key2[0]), .B1(
        Key2[64]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1871) );
  MUX2_X1 Midori_rounds_U253 ( .A(Midori_rounds_n1360), .B(
        Midori_rounds_SR_Result1[9]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[9]) );
  XNOR2_X1 Midori_rounds_U252 ( .A(Midori_rounds_SR_Result1[9]), .B(
        Midori_rounds_n1997), .ZN(Midori_rounds_n1360) );
  AOI22_X1 Midori_rounds_U251 ( .A1(Midori_rounds_n1269), .A2(Key1[9]), .B1(
        Key1[73]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1997) );
  MUX2_X1 Midori_rounds_U250 ( .A(Midori_rounds_n1359), .B(
        Midori_rounds_SR_Result1[8]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[8]) );
  XNOR2_X1 Midori_rounds_U249 ( .A(Midori_rounds_SR_Result1[8]), .B(
        Midori_rounds_n2057), .ZN(Midori_rounds_n1359) );
  XOR2_X1 Midori_rounds_U248 ( .A(Midori_rounds_round_Constant[2]), .B(
        Midori_rounds_n1358), .Z(Midori_rounds_n2057) );
  AOI22_X1 Midori_rounds_U247 ( .A1(Midori_rounds_n1269), .A2(Key1[8]), .B1(
        Key1[72]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1358) );
  MUX2_X1 Midori_rounds_U246 ( .A(Midori_rounds_n1357), .B(
        Midori_rounds_SR_Result1[7]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[7]) );
  XNOR2_X1 Midori_rounds_U245 ( .A(Midori_rounds_SR_Result1[47]), .B(
        Midori_rounds_n2000), .ZN(Midori_rounds_n1357) );
  AOI22_X1 Midori_rounds_U244 ( .A1(Midori_rounds_n1269), .A2(Key1[7]), .B1(
        Key1[71]), .B2(Midori_rounds_n1275), .ZN(Midori_rounds_n2000) );
  MUX2_X1 Midori_rounds_U243 ( .A(Midori_rounds_n1356), .B(
        Midori_rounds_SR_Result1[6]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[6]) );
  XNOR2_X1 Midori_rounds_U242 ( .A(Midori_rounds_SR_Result1[46]), .B(
        Midori_rounds_n2003), .ZN(Midori_rounds_n1356) );
  AOI22_X1 Midori_rounds_U241 ( .A1(Midori_rounds_n1269), .A2(Key1[6]), .B1(
        Key1[70]), .B2(Midori_rounds_n1275), .ZN(Midori_rounds_n2003) );
  MUX2_X1 Midori_rounds_U240 ( .A(Midori_rounds_n1355), .B(
        Midori_rounds_SR_Result1[63]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[63]) );
  XNOR2_X1 Midori_rounds_U239 ( .A(Midori_rounds_SR_Result1[63]), .B(
        Midori_rounds_n1874), .ZN(Midori_rounds_n1355) );
  AOI22_X1 Midori_rounds_U238 ( .A1(Midori_rounds_n1269), .A2(Key1[63]), .B1(
        Key1[127]), .B2(Midori_rounds_n1275), .ZN(Midori_rounds_n1874) );
  MUX2_X1 Midori_rounds_U237 ( .A(Midori_rounds_n1354), .B(
        Midori_rounds_SR_Result1[62]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[62]) );
  XNOR2_X1 Midori_rounds_U236 ( .A(Midori_rounds_SR_Result1[62]), .B(
        Midori_rounds_n1877), .ZN(Midori_rounds_n1354) );
  AOI22_X1 Midori_rounds_U235 ( .A1(Midori_rounds_n1269), .A2(Key1[62]), .B1(
        Key1[126]), .B2(Midori_rounds_n1275), .ZN(Midori_rounds_n1877) );
  MUX2_X1 Midori_rounds_U234 ( .A(Midori_rounds_n1353), .B(
        Midori_rounds_SR_Result1[61]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[61]) );
  XNOR2_X1 Midori_rounds_U233 ( .A(Midori_rounds_SR_Result1[61]), .B(
        Midori_rounds_n1880), .ZN(Midori_rounds_n1353) );
  AOI22_X1 Midori_rounds_U232 ( .A1(Midori_rounds_n1269), .A2(Key1[61]), .B1(
        Key1[125]), .B2(Midori_rounds_n1275), .ZN(Midori_rounds_n1880) );
  MUX2_X1 Midori_rounds_U231 ( .A(Midori_rounds_n1352), .B(
        Midori_rounds_SR_Result1[60]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[60]) );
  XNOR2_X1 Midori_rounds_U230 ( .A(Midori_rounds_SR_Result1[60]), .B(
        Midori_rounds_n2018), .ZN(Midori_rounds_n1352) );
  XOR2_X1 Midori_rounds_U229 ( .A(Midori_rounds_round_Constant[15]), .B(
        Midori_rounds_n1351), .Z(Midori_rounds_n2018) );
  AOI22_X1 Midori_rounds_U228 ( .A1(Midori_rounds_n1269), .A2(Key1[60]), .B1(
        Key1[124]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1351) );
  MUX2_X1 Midori_rounds_U227 ( .A(Midori_rounds_n1350), .B(
        Midori_rounds_SR_Result1[5]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[5]) );
  XNOR2_X1 Midori_rounds_U226 ( .A(Midori_rounds_SR_Result1[45]), .B(
        Midori_rounds_n2006), .ZN(Midori_rounds_n1350) );
  AOI22_X1 Midori_rounds_U225 ( .A1(Midori_rounds_n1269), .A2(Key1[5]), .B1(
        Key1[69]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n2006) );
  MUX2_X1 Midori_rounds_U224 ( .A(Midori_rounds_n1349), .B(
        Midori_rounds_SR_Result1[59]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[59]) );
  XNOR2_X1 Midori_rounds_U223 ( .A(Midori_rounds_SR_Result1[35]), .B(
        Midori_rounds_n1883), .ZN(Midori_rounds_n1349) );
  AOI22_X1 Midori_rounds_U222 ( .A1(Midori_rounds_n1269), .A2(Key1[59]), .B1(
        Key1[123]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1883) );
  MUX2_X1 Midori_rounds_U221 ( .A(Midori_rounds_n1348), .B(
        Midori_rounds_SR_Result1[58]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[58]) );
  XNOR2_X1 Midori_rounds_U220 ( .A(Midori_rounds_SR_Result1[34]), .B(
        Midori_rounds_n1886), .ZN(Midori_rounds_n1348) );
  AOI22_X1 Midori_rounds_U219 ( .A1(Midori_rounds_n1269), .A2(Key1[58]), .B1(
        Key1[122]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1886) );
  MUX2_X1 Midori_rounds_U218 ( .A(Midori_rounds_n1347), .B(
        Midori_rounds_SR_Result1[57]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[57]) );
  XNOR2_X1 Midori_rounds_U217 ( .A(Midori_rounds_SR_Result1[33]), .B(
        Midori_rounds_n1889), .ZN(Midori_rounds_n1347) );
  AOI22_X1 Midori_rounds_U216 ( .A1(Midori_rounds_n1269), .A2(Key1[57]), .B1(
        Key1[121]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1889) );
  MUX2_X1 Midori_rounds_U215 ( .A(Midori_rounds_n1346), .B(
        Midori_rounds_SR_Result1[56]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[56]) );
  XNOR2_X1 Midori_rounds_U214 ( .A(Midori_rounds_SR_Result1[32]), .B(
        Midori_rounds_n2021), .ZN(Midori_rounds_n1346) );
  XOR2_X1 Midori_rounds_U213 ( .A(Midori_rounds_round_Constant[14]), .B(
        Midori_rounds_n1345), .Z(Midori_rounds_n2021) );
  AOI22_X1 Midori_rounds_U212 ( .A1(Midori_rounds_n1269), .A2(Key1[56]), .B1(
        Key1[120]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1345) );
  MUX2_X1 Midori_rounds_U211 ( .A(Midori_rounds_n1344), .B(
        Midori_rounds_SR_Result1[55]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[55]) );
  XNOR2_X1 Midori_rounds_U210 ( .A(Midori_rounds_SR_Result1[7]), .B(
        Midori_rounds_n1892), .ZN(Midori_rounds_n1344) );
  AOI22_X1 Midori_rounds_U209 ( .A1(Midori_rounds_n1268), .A2(Key1[55]), .B1(
        Key1[119]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1892) );
  MUX2_X1 Midori_rounds_U208 ( .A(Midori_rounds_n1343), .B(
        Midori_rounds_SR_Result1[54]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[54]) );
  XNOR2_X1 Midori_rounds_U207 ( .A(Midori_rounds_SR_Result1[6]), .B(
        Midori_rounds_n1895), .ZN(Midori_rounds_n1343) );
  AOI22_X1 Midori_rounds_U206 ( .A1(Midori_rounds_n1268), .A2(Key1[54]), .B1(
        Key1[118]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1895) );
  MUX2_X1 Midori_rounds_U205 ( .A(Midori_rounds_n1342), .B(
        Midori_rounds_SR_Result1[53]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[53]) );
  XNOR2_X1 Midori_rounds_U204 ( .A(Midori_rounds_SR_Result1[5]), .B(
        Midori_rounds_n1898), .ZN(Midori_rounds_n1342) );
  AOI22_X1 Midori_rounds_U203 ( .A1(Midori_rounds_n1268), .A2(Key1[53]), .B1(
        Key1[117]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1898) );
  MUX2_X1 Midori_rounds_U202 ( .A(Midori_rounds_n1341), .B(
        Midori_rounds_SR_Result1[52]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[52]) );
  XNOR2_X1 Midori_rounds_U201 ( .A(Midori_rounds_SR_Result1[4]), .B(
        Midori_rounds_n2024), .ZN(Midori_rounds_n1341) );
  XOR2_X1 Midori_rounds_U200 ( .A(Midori_rounds_round_Constant[13]), .B(
        Midori_rounds_n1340), .Z(Midori_rounds_n2024) );
  AOI22_X1 Midori_rounds_U199 ( .A1(Midori_rounds_n1268), .A2(Key1[52]), .B1(
        Key1[116]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1340) );
  MUX2_X1 Midori_rounds_U198 ( .A(Midori_rounds_n1339), .B(
        Midori_rounds_SR_Result1[51]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[51]) );
  XNOR2_X1 Midori_rounds_U197 ( .A(Midori_rounds_SR_Result1[27]), .B(
        Midori_rounds_n1901), .ZN(Midori_rounds_n1339) );
  AOI22_X1 Midori_rounds_U196 ( .A1(Midori_rounds_n1268), .A2(Key1[51]), .B1(
        Key1[115]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1901) );
  MUX2_X1 Midori_rounds_U195 ( .A(Midori_rounds_n1338), .B(
        Midori_rounds_SR_Result1[50]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[50]) );
  XNOR2_X1 Midori_rounds_U194 ( .A(Midori_rounds_SR_Result1[26]), .B(
        Midori_rounds_n1904), .ZN(Midori_rounds_n1338) );
  AOI22_X1 Midori_rounds_U193 ( .A1(Midori_rounds_n1268), .A2(Key1[50]), .B1(
        Key1[114]), .B2(Midori_rounds_n1279), .ZN(Midori_rounds_n1904) );
  MUX2_X1 Midori_rounds_U192 ( .A(Midori_rounds_n1337), .B(
        Midori_rounds_SR_Result1[4]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[4]) );
  XNOR2_X1 Midori_rounds_U191 ( .A(Midori_rounds_SR_Result1[44]), .B(
        Midori_rounds_n2060), .ZN(Midori_rounds_n1337) );
  XOR2_X1 Midori_rounds_U190 ( .A(Midori_rounds_round_Constant[1]), .B(
        Midori_rounds_n1336), .Z(Midori_rounds_n2060) );
  AOI22_X1 Midori_rounds_U189 ( .A1(Midori_rounds_n1268), .A2(Key1[4]), .B1(
        Key1[68]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1336) );
  MUX2_X1 Midori_rounds_U188 ( .A(Midori_rounds_n1335), .B(
        Midori_rounds_SR_Result1[49]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[49]) );
  XNOR2_X1 Midori_rounds_U187 ( .A(Midori_rounds_SR_Result1[25]), .B(
        Midori_rounds_n1907), .ZN(Midori_rounds_n1335) );
  AOI22_X1 Midori_rounds_U186 ( .A1(Midori_rounds_n1268), .A2(Key1[49]), .B1(
        Key1[113]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1907) );
  MUX2_X1 Midori_rounds_U185 ( .A(Midori_rounds_n1334), .B(
        Midori_rounds_SR_Result1[48]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[48]) );
  XNOR2_X1 Midori_rounds_U184 ( .A(Midori_rounds_SR_Result1[24]), .B(
        Midori_rounds_n2027), .ZN(Midori_rounds_n1334) );
  XOR2_X1 Midori_rounds_U183 ( .A(Midori_rounds_round_Constant[12]), .B(
        Midori_rounds_n1333), .Z(Midori_rounds_n2027) );
  AOI22_X1 Midori_rounds_U182 ( .A1(Midori_rounds_n1268), .A2(Key1[48]), .B1(
        Key1[112]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1333) );
  MUX2_X1 Midori_rounds_U181 ( .A(Midori_rounds_n1332), .B(
        Midori_rounds_SR_Result1[47]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[47]) );
  XNOR2_X1 Midori_rounds_U180 ( .A(Midori_rounds_SR_Result1[43]), .B(
        Midori_rounds_n1910), .ZN(Midori_rounds_n1332) );
  AOI22_X1 Midori_rounds_U179 ( .A1(Midori_rounds_n1268), .A2(Key1[47]), .B1(
        Key1[111]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1910) );
  MUX2_X1 Midori_rounds_U178 ( .A(Midori_rounds_n1331), .B(
        Midori_rounds_SR_Result1[46]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[46]) );
  XNOR2_X1 Midori_rounds_U177 ( .A(Midori_rounds_SR_Result1[42]), .B(
        Midori_rounds_n1913), .ZN(Midori_rounds_n1331) );
  AOI22_X1 Midori_rounds_U176 ( .A1(Midori_rounds_n1268), .A2(Key1[46]), .B1(
        Key1[110]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1913) );
  MUX2_X1 Midori_rounds_U175 ( .A(Midori_rounds_n1330), .B(
        Midori_rounds_SR_Result1[45]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[45]) );
  XNOR2_X1 Midori_rounds_U174 ( .A(Midori_rounds_SR_Result1[41]), .B(
        Midori_rounds_n1916), .ZN(Midori_rounds_n1330) );
  AOI22_X1 Midori_rounds_U173 ( .A1(Midori_rounds_n1268), .A2(Key1[45]), .B1(
        Key1[109]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1916) );
  MUX2_X1 Midori_rounds_U172 ( .A(Midori_rounds_n1329), .B(
        Midori_rounds_SR_Result1[44]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[44]) );
  XNOR2_X1 Midori_rounds_U171 ( .A(Midori_rounds_SR_Result1[40]), .B(
        Midori_rounds_n2030), .ZN(Midori_rounds_n1329) );
  XOR2_X1 Midori_rounds_U170 ( .A(Midori_rounds_round_Constant[11]), .B(
        Midori_rounds_n1328), .Z(Midori_rounds_n2030) );
  AOI22_X1 Midori_rounds_U169 ( .A1(Midori_rounds_n1268), .A2(Key1[44]), .B1(
        Key1[108]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1328) );
  MUX2_X1 Midori_rounds_U168 ( .A(Midori_rounds_n1327), .B(
        Midori_rounds_SR_Result1[43]), .S(Midori_rounds_n1243), .Z(
        Midori_rounds_mul_input1[43]) );
  XNOR2_X1 Midori_rounds_U167 ( .A(Midori_rounds_SR_Result1[55]), .B(
        Midori_rounds_n1919), .ZN(Midori_rounds_n1327) );
  AOI22_X1 Midori_rounds_U166 ( .A1(round_Signal[0]), .A2(Key1[43]), .B1(
        Key1[107]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1919) );
  MUX2_X1 Midori_rounds_U165 ( .A(Midori_rounds_n1326), .B(
        Midori_rounds_SR_Result1[42]), .S(Midori_rounds_n1249), .Z(
        Midori_rounds_mul_input1[42]) );
  XNOR2_X1 Midori_rounds_U164 ( .A(Midori_rounds_SR_Result1[54]), .B(
        Midori_rounds_n1922), .ZN(Midori_rounds_n1326) );
  AOI22_X1 Midori_rounds_U163 ( .A1(round_Signal[0]), .A2(Key1[42]), .B1(
        Key1[106]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1922) );
  MUX2_X1 Midori_rounds_U162 ( .A(Midori_rounds_n1325), .B(
        Midori_rounds_SR_Result1[41]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[41]) );
  XNOR2_X1 Midori_rounds_U161 ( .A(Midori_rounds_SR_Result1[53]), .B(
        Midori_rounds_n1925), .ZN(Midori_rounds_n1325) );
  AOI22_X1 Midori_rounds_U160 ( .A1(Midori_rounds_n1267), .A2(Key1[41]), .B1(
        Key1[105]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1925) );
  MUX2_X1 Midori_rounds_U159 ( .A(Midori_rounds_n1324), .B(
        Midori_rounds_SR_Result1[40]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[40]) );
  XNOR2_X1 Midori_rounds_U158 ( .A(Midori_rounds_SR_Result1[52]), .B(
        Midori_rounds_n2033), .ZN(Midori_rounds_n1324) );
  XOR2_X1 Midori_rounds_U157 ( .A(Midori_rounds_round_Constant[10]), .B(
        Midori_rounds_n1323), .Z(Midori_rounds_n2033) );
  AOI22_X1 Midori_rounds_U156 ( .A1(round_Signal[0]), .A2(Key1[40]), .B1(
        Key1[104]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1323) );
  MUX2_X1 Midori_rounds_U155 ( .A(Midori_rounds_n1322), .B(
        Midori_rounds_SR_Result1[3]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[3]) );
  XNOR2_X1 Midori_rounds_U154 ( .A(Midori_rounds_SR_Result1[51]), .B(
        Midori_rounds_n2009), .ZN(Midori_rounds_n1322) );
  AOI22_X1 Midori_rounds_U153 ( .A1(Midori_rounds_n1267), .A2(Key1[3]), .B1(
        Key1[67]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n2009) );
  MUX2_X1 Midori_rounds_U152 ( .A(Midori_rounds_n1321), .B(
        Midori_rounds_SR_Result1[39]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[39]) );
  XNOR2_X1 Midori_rounds_U151 ( .A(Midori_rounds_SR_Result1[19]), .B(
        Midori_rounds_n1928), .ZN(Midori_rounds_n1321) );
  AOI22_X1 Midori_rounds_U150 ( .A1(round_Signal[0]), .A2(Key1[39]), .B1(
        Key1[103]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1928) );
  MUX2_X1 Midori_rounds_U149 ( .A(Midori_rounds_n1320), .B(
        Midori_rounds_SR_Result1[38]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[38]) );
  XNOR2_X1 Midori_rounds_U148 ( .A(Midori_rounds_SR_Result1[18]), .B(
        Midori_rounds_n1931), .ZN(Midori_rounds_n1320) );
  AOI22_X1 Midori_rounds_U147 ( .A1(round_Signal[0]), .A2(Key1[38]), .B1(
        Key1[102]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1931) );
  MUX2_X1 Midori_rounds_U146 ( .A(Midori_rounds_n1319), .B(
        Midori_rounds_SR_Result1[37]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[37]) );
  XNOR2_X1 Midori_rounds_U145 ( .A(Midori_rounds_SR_Result1[17]), .B(
        Midori_rounds_n1934), .ZN(Midori_rounds_n1319) );
  AOI22_X1 Midori_rounds_U144 ( .A1(round_Signal[0]), .A2(Key1[37]), .B1(
        Key1[101]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1934) );
  MUX2_X1 Midori_rounds_U143 ( .A(Midori_rounds_n1318), .B(
        Midori_rounds_SR_Result1[36]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[36]) );
  XNOR2_X1 Midori_rounds_U142 ( .A(Midori_rounds_SR_Result1[16]), .B(
        Midori_rounds_n2036), .ZN(Midori_rounds_n1318) );
  XOR2_X1 Midori_rounds_U141 ( .A(Midori_rounds_round_Constant[9]), .B(
        Midori_rounds_n1317), .Z(Midori_rounds_n2036) );
  AOI22_X1 Midori_rounds_U140 ( .A1(round_Signal[0]), .A2(Key1[36]), .B1(
        Key1[100]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1317) );
  MUX2_X1 Midori_rounds_U139 ( .A(Midori_rounds_n1316), .B(
        Midori_rounds_SR_Result1[35]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[35]) );
  XNOR2_X1 Midori_rounds_U138 ( .A(Midori_rounds_SR_Result1[15]), .B(
        Midori_rounds_n1937), .ZN(Midori_rounds_n1316) );
  AOI22_X1 Midori_rounds_U137 ( .A1(round_Signal[0]), .A2(Key1[35]), .B1(
        Key1[99]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1937) );
  MUX2_X1 Midori_rounds_U136 ( .A(Midori_rounds_n1315), .B(
        Midori_rounds_SR_Result1[34]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[34]) );
  XNOR2_X1 Midori_rounds_U135 ( .A(Midori_rounds_SR_Result1[14]), .B(
        Midori_rounds_n1940), .ZN(Midori_rounds_n1315) );
  AOI22_X1 Midori_rounds_U134 ( .A1(round_Signal[0]), .A2(Key1[34]), .B1(
        Key1[98]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1940) );
  MUX2_X1 Midori_rounds_U133 ( .A(Midori_rounds_n1314), .B(
        Midori_rounds_SR_Result1[33]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[33]) );
  XNOR2_X1 Midori_rounds_U132 ( .A(Midori_rounds_SR_Result1[13]), .B(
        Midori_rounds_n1943), .ZN(Midori_rounds_n1314) );
  AOI22_X1 Midori_rounds_U131 ( .A1(Midori_rounds_n1267), .A2(Key1[33]), .B1(
        Key1[97]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1943) );
  MUX2_X1 Midori_rounds_U130 ( .A(Midori_rounds_n1313), .B(
        Midori_rounds_SR_Result1[32]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[32]) );
  XNOR2_X1 Midori_rounds_U129 ( .A(Midori_rounds_SR_Result1[12]), .B(
        Midori_rounds_n2039), .ZN(Midori_rounds_n1313) );
  XOR2_X1 Midori_rounds_U128 ( .A(Midori_rounds_round_Constant[8]), .B(
        Midori_rounds_n1312), .Z(Midori_rounds_n2039) );
  AOI22_X1 Midori_rounds_U127 ( .A1(Midori_rounds_n1267), .A2(Key1[32]), .B1(
        Key1[96]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1312) );
  MUX2_X1 Midori_rounds_U126 ( .A(Midori_rounds_n1311), .B(
        Midori_rounds_SR_Result1[31]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[31]) );
  XNOR2_X1 Midori_rounds_U125 ( .A(Midori_rounds_SR_Result1[3]), .B(
        Midori_rounds_n1946), .ZN(Midori_rounds_n1311) );
  AOI22_X1 Midori_rounds_U124 ( .A1(Midori_rounds_n1267), .A2(Key1[31]), .B1(
        Key1[95]), .B2(Midori_rounds_n1281), .ZN(Midori_rounds_n1946) );
  MUX2_X1 Midori_rounds_U123 ( .A(Midori_rounds_n1310), .B(
        Midori_rounds_SR_Result1[30]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[30]) );
  XNOR2_X1 Midori_rounds_U122 ( .A(Midori_rounds_SR_Result1[2]), .B(
        Midori_rounds_n1949), .ZN(Midori_rounds_n1310) );
  AOI22_X1 Midori_rounds_U121 ( .A1(round_Signal[0]), .A2(Key1[30]), .B1(
        Key1[94]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1949) );
  MUX2_X1 Midori_rounds_U120 ( .A(Midori_rounds_n1309), .B(
        Midori_rounds_SR_Result1[2]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[2]) );
  XNOR2_X1 Midori_rounds_U119 ( .A(Midori_rounds_SR_Result1[50]), .B(
        Midori_rounds_n2012), .ZN(Midori_rounds_n1309) );
  AOI22_X1 Midori_rounds_U118 ( .A1(round_Signal[0]), .A2(Key1[2]), .B1(
        Key1[66]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n2012) );
  MUX2_X1 Midori_rounds_U117 ( .A(Midori_rounds_n1308), .B(
        Midori_rounds_SR_Result1[29]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[29]) );
  XNOR2_X1 Midori_rounds_U116 ( .A(Midori_rounds_SR_Result1[1]), .B(
        Midori_rounds_n1952), .ZN(Midori_rounds_n1308) );
  AOI22_X1 Midori_rounds_U115 ( .A1(Midori_rounds_n1267), .A2(Key1[29]), .B1(
        Key1[93]), .B2(Midori_rounds_n1278), .ZN(Midori_rounds_n1952) );
  MUX2_X1 Midori_rounds_U114 ( .A(Midori_rounds_n1307), .B(
        Midori_rounds_SR_Result1[28]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[28]) );
  XNOR2_X1 Midori_rounds_U113 ( .A(Midori_rounds_SR_Result1[0]), .B(
        Midori_rounds_n2042), .ZN(Midori_rounds_n1307) );
  XOR2_X1 Midori_rounds_U112 ( .A(Midori_rounds_round_Constant[7]), .B(
        Midori_rounds_n1306), .Z(Midori_rounds_n2042) );
  AOI22_X1 Midori_rounds_U111 ( .A1(round_Signal[0]), .A2(Key1[28]), .B1(
        Key1[92]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1306) );
  MUX2_X1 Midori_rounds_U110 ( .A(Midori_rounds_n1305), .B(
        Midori_rounds_SR_Result1[27]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[27]) );
  XNOR2_X1 Midori_rounds_U109 ( .A(Midori_rounds_SR_Result1[31]), .B(
        Midori_rounds_n1955), .ZN(Midori_rounds_n1305) );
  AOI22_X1 Midori_rounds_U108 ( .A1(round_Signal[0]), .A2(Key1[27]), .B1(
        Key1[91]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1955) );
  MUX2_X1 Midori_rounds_U107 ( .A(Midori_rounds_n1304), .B(
        Midori_rounds_SR_Result1[26]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[26]) );
  XNOR2_X1 Midori_rounds_U106 ( .A(Midori_rounds_SR_Result1[30]), .B(
        Midori_rounds_n1958), .ZN(Midori_rounds_n1304) );
  AOI22_X1 Midori_rounds_U105 ( .A1(round_Signal[0]), .A2(Key1[26]), .B1(
        Key1[90]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1958) );
  MUX2_X1 Midori_rounds_U104 ( .A(Midori_rounds_n1303), .B(
        Midori_rounds_SR_Result1[25]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[25]) );
  XNOR2_X1 Midori_rounds_U103 ( .A(Midori_rounds_SR_Result1[29]), .B(
        Midori_rounds_n1961), .ZN(Midori_rounds_n1303) );
  AOI22_X1 Midori_rounds_U102 ( .A1(Midori_rounds_n1267), .A2(Key1[25]), .B1(
        Key1[89]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1961) );
  MUX2_X1 Midori_rounds_U101 ( .A(Midori_rounds_n1302), .B(
        Midori_rounds_SR_Result1[24]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[24]) );
  XNOR2_X1 Midori_rounds_U100 ( .A(Midori_rounds_SR_Result1[28]), .B(
        Midori_rounds_n2045), .ZN(Midori_rounds_n1302) );
  XOR2_X1 Midori_rounds_U99 ( .A(Midori_rounds_round_Constant[6]), .B(
        Midori_rounds_n1301), .Z(Midori_rounds_n2045) );
  AOI22_X1 Midori_rounds_U98 ( .A1(Midori_rounds_n1267), .A2(Key1[24]), .B1(
        Key1[88]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1301) );
  MUX2_X1 Midori_rounds_U97 ( .A(Midori_rounds_n1300), .B(
        Midori_rounds_SR_Result1[23]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[23]) );
  XNOR2_X1 Midori_rounds_U96 ( .A(Midori_rounds_SR_Result1[59]), .B(
        Midori_rounds_n1964), .ZN(Midori_rounds_n1300) );
  AOI22_X1 Midori_rounds_U95 ( .A1(round_Signal[0]), .A2(Key1[23]), .B1(
        Key1[87]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1964) );
  MUX2_X1 Midori_rounds_U94 ( .A(Midori_rounds_n1299), .B(
        Midori_rounds_SR_Result1[22]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[22]) );
  XNOR2_X1 Midori_rounds_U93 ( .A(Midori_rounds_SR_Result1[58]), .B(
        Midori_rounds_n1967), .ZN(Midori_rounds_n1299) );
  AOI22_X1 Midori_rounds_U92 ( .A1(round_Signal[0]), .A2(Key1[22]), .B1(
        Key1[86]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1967) );
  MUX2_X1 Midori_rounds_U91 ( .A(Midori_rounds_n1298), .B(
        Midori_rounds_SR_Result1[21]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[21]) );
  XNOR2_X1 Midori_rounds_U90 ( .A(Midori_rounds_SR_Result1[57]), .B(
        Midori_rounds_n1970), .ZN(Midori_rounds_n1298) );
  AOI22_X1 Midori_rounds_U89 ( .A1(Midori_rounds_n1267), .A2(Key1[21]), .B1(
        Key1[85]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1970) );
  MUX2_X1 Midori_rounds_U88 ( .A(Midori_rounds_n1297), .B(
        Midori_rounds_SR_Result1[20]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[20]) );
  XNOR2_X1 Midori_rounds_U87 ( .A(Midori_rounds_SR_Result1[56]), .B(
        Midori_rounds_n2048), .ZN(Midori_rounds_n1297) );
  MUX2_X1 Midori_rounds_U86 ( .A(Midori_rounds_n1296), .B(
        Midori_rounds_SR_Result1[1]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[1]) );
  XNOR2_X1 Midori_rounds_U85 ( .A(Midori_rounds_SR_Result1[49]), .B(
        Midori_rounds_n2015), .ZN(Midori_rounds_n1296) );
  AOI22_X1 Midori_rounds_U84 ( .A1(Midori_rounds_n1267), .A2(Key1[1]), .B1(
        Key1[65]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n2015) );
  MUX2_X1 Midori_rounds_U83 ( .A(Midori_rounds_n1295), .B(
        Midori_rounds_SR_Result1[19]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[19]) );
  XNOR2_X1 Midori_rounds_U82 ( .A(Midori_rounds_SR_Result1[39]), .B(
        Midori_rounds_n1973), .ZN(Midori_rounds_n1295) );
  AOI22_X1 Midori_rounds_U81 ( .A1(Midori_rounds_n1267), .A2(Key1[19]), .B1(
        Key1[83]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1973) );
  MUX2_X1 Midori_rounds_U80 ( .A(Midori_rounds_n1294), .B(
        Midori_rounds_SR_Result1[18]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[18]) );
  XNOR2_X1 Midori_rounds_U79 ( .A(Midori_rounds_SR_Result1[38]), .B(
        Midori_rounds_n1976), .ZN(Midori_rounds_n1294) );
  AOI22_X1 Midori_rounds_U78 ( .A1(Midori_rounds_n1267), .A2(Key1[18]), .B1(
        Key1[82]), .B2(Midori_rounds_n1277), .ZN(Midori_rounds_n1976) );
  MUX2_X1 Midori_rounds_U77 ( .A(Midori_rounds_n1293), .B(
        Midori_rounds_SR_Result1[17]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[17]) );
  XNOR2_X1 Midori_rounds_U76 ( .A(Midori_rounds_SR_Result1[37]), .B(
        Midori_rounds_n1979), .ZN(Midori_rounds_n1293) );
  AOI22_X1 Midori_rounds_U75 ( .A1(Midori_rounds_n1267), .A2(Key1[17]), .B1(
        Key1[81]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1979) );
  MUX2_X1 Midori_rounds_U74 ( .A(Midori_rounds_n1292), .B(
        Midori_rounds_SR_Result1[16]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[16]) );
  XNOR2_X1 Midori_rounds_U73 ( .A(Midori_rounds_SR_Result1[36]), .B(
        Midori_rounds_n2051), .ZN(Midori_rounds_n1292) );
  XOR2_X1 Midori_rounds_U72 ( .A(Midori_rounds_round_Constant[4]), .B(
        Midori_rounds_n1291), .Z(Midori_rounds_n2051) );
  AOI22_X1 Midori_rounds_U71 ( .A1(Midori_rounds_n1267), .A2(Key1[16]), .B1(
        Key1[80]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1291) );
  MUX2_X1 Midori_rounds_U70 ( .A(Midori_rounds_n1290), .B(
        Midori_rounds_SR_Result1[15]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[15]) );
  XNOR2_X1 Midori_rounds_U69 ( .A(Midori_rounds_SR_Result1[23]), .B(
        Midori_rounds_n1982), .ZN(Midori_rounds_n1290) );
  AOI22_X1 Midori_rounds_U68 ( .A1(Midori_rounds_n1267), .A2(Key1[15]), .B1(
        Key1[79]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1982) );
  MUX2_X1 Midori_rounds_U67 ( .A(Midori_rounds_n1289), .B(
        Midori_rounds_SR_Result1[14]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[14]) );
  XNOR2_X1 Midori_rounds_U66 ( .A(Midori_rounds_SR_Result1[22]), .B(
        Midori_rounds_n1985), .ZN(Midori_rounds_n1289) );
  AOI22_X1 Midori_rounds_U65 ( .A1(Midori_rounds_n1267), .A2(Key1[14]), .B1(
        Key1[78]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1985) );
  MUX2_X1 Midori_rounds_U64 ( .A(Midori_rounds_n1288), .B(
        Midori_rounds_SR_Result1[13]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[13]) );
  XNOR2_X1 Midori_rounds_U63 ( .A(Midori_rounds_SR_Result1[21]), .B(
        Midori_rounds_n1988), .ZN(Midori_rounds_n1288) );
  AOI22_X1 Midori_rounds_U62 ( .A1(Midori_rounds_n1267), .A2(Key1[13]), .B1(
        Key1[77]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1988) );
  MUX2_X1 Midori_rounds_U61 ( .A(Midori_rounds_n1287), .B(
        Midori_rounds_SR_Result1[12]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[12]) );
  XNOR2_X1 Midori_rounds_U60 ( .A(Midori_rounds_SR_Result1[20]), .B(
        Midori_rounds_n2054), .ZN(Midori_rounds_n1287) );
  XOR2_X1 Midori_rounds_U59 ( .A(Midori_rounds_round_Constant[3]), .B(
        Midori_rounds_n1286), .Z(Midori_rounds_n2054) );
  AOI22_X1 Midori_rounds_U58 ( .A1(Midori_rounds_n1267), .A2(Key1[12]), .B1(
        Key1[76]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1286) );
  MUX2_X1 Midori_rounds_U57 ( .A(Midori_rounds_n1285), .B(
        Midori_rounds_SR_Result1[11]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[11]) );
  XNOR2_X1 Midori_rounds_U56 ( .A(Midori_rounds_SR_Result1[11]), .B(
        Midori_rounds_n1991), .ZN(Midori_rounds_n1285) );
  AOI22_X1 Midori_rounds_U55 ( .A1(Midori_rounds_n1267), .A2(Key1[11]), .B1(
        Key1[75]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1991) );
  MUX2_X1 Midori_rounds_U54 ( .A(Midori_rounds_n1284), .B(
        Midori_rounds_SR_Result1[10]), .S(Midori_rounds_n1242), .Z(
        Midori_rounds_mul_input1[10]) );
  XNOR2_X1 Midori_rounds_U53 ( .A(Midori_rounds_SR_Result1[10]), .B(
        Midori_rounds_n1994), .ZN(Midori_rounds_n1284) );
  AOI22_X1 Midori_rounds_U52 ( .A1(Midori_rounds_n1267), .A2(Key1[10]), .B1(
        Key1[74]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1994) );
  MUX2_X1 Midori_rounds_U51 ( .A(Midori_rounds_n1283), .B(
        Midori_rounds_SR_Result1[0]), .S(Midori_rounds_n1248), .Z(
        Midori_rounds_mul_input1[0]) );
  XNOR2_X1 Midori_rounds_U50 ( .A(Midori_rounds_SR_Result1[48]), .B(
        Midori_rounds_n2063), .ZN(Midori_rounds_n1283) );
  XOR2_X1 Midori_rounds_U49 ( .A(Midori_rounds_round_Constant[0]), .B(
        Midori_rounds_n1282), .Z(Midori_rounds_n2063) );
  AOI22_X1 Midori_rounds_U48 ( .A1(Midori_rounds_n1267), .A2(Key1[0]), .B1(
        Key1[64]), .B2(Midori_rounds_n1276), .ZN(Midori_rounds_n1282) );
  INV_X1 Midori_rounds_U47 ( .A(Midori_rounds_n1275), .ZN(Midori_rounds_n1268)
         );
  BUF_X1 Midori_rounds_U46 ( .A(Midori_rounds_n1275), .Z(Midori_rounds_n1279)
         );
  INV_X1 Midori_rounds_U45 ( .A(enc_dec), .ZN(Midori_rounds_n1490) );
  BUF_X1 Midori_rounds_U44 ( .A(Midori_rounds_n1490), .Z(Midori_rounds_n1247)
         );
  BUF_X1 Midori_rounds_U43 ( .A(Midori_rounds_n1247), .Z(Midori_rounds_n1243)
         );
  INV_X1 Midori_rounds_U42 ( .A(Midori_rounds_n1275), .ZN(Midori_rounds_n1269)
         );
  BUF_X2 Midori_rounds_U41 ( .A(Midori_rounds_n2066), .Z(Midori_rounds_n1265)
         );
  BUF_X1 Midori_rounds_U40 ( .A(Midori_rounds_n1490), .Z(Midori_rounds_n1246)
         );
  NOR2_X1 Midori_rounds_U39 ( .A1(reset), .A2(Midori_rounds_n1246), .ZN(
        Midori_rounds_n2064) );
  BUF_X1 Midori_rounds_U38 ( .A(Midori_rounds_n1247), .Z(Midori_rounds_n1242)
         );
  BUF_X1 Midori_rounds_U37 ( .A(Midori_rounds_n2066), .Z(Midori_rounds_n1262)
         );
  BUF_X1 Midori_rounds_U36 ( .A(Midori_rounds_n2064), .Z(Midori_rounds_n1255)
         );
  BUF_X1 Midori_rounds_U35 ( .A(Midori_rounds_n1242), .Z(Midori_rounds_n1248)
         );
  BUF_X1 Midori_rounds_U34 ( .A(Midori_rounds_n1243), .Z(Midori_rounds_n1249)
         );
  BUF_X1 Midori_rounds_U33 ( .A(Midori_rounds_n2064), .Z(Midori_rounds_n1257)
         );
  BUF_X1 Midori_rounds_U32 ( .A(Midori_rounds_n1257), .Z(Midori_rounds_n1251)
         );
  BUF_X1 Midori_rounds_U31 ( .A(Midori_rounds_n2066), .Z(Midori_rounds_n1266)
         );
  BUF_X1 Midori_rounds_U30 ( .A(Midori_rounds_n1257), .Z(Midori_rounds_n1253)
         );
  BUF_X1 Midori_rounds_U29 ( .A(Midori_rounds_n2066), .Z(Midori_rounds_n1264)
         );
  BUF_X1 Midori_rounds_U28 ( .A(Midori_rounds_n2064), .Z(Midori_rounds_n1256)
         );
  BUF_X1 Midori_rounds_U27 ( .A(Midori_rounds_n1256), .Z(Midori_rounds_n1259)
         );
  BUF_X1 Midori_rounds_U26 ( .A(Midori_rounds_n2066), .Z(Midori_rounds_n1263)
         );
  BUF_X1 Midori_rounds_U25 ( .A(Midori_rounds_n2064), .Z(Midori_rounds_n1258)
         );
  BUF_X1 Midori_rounds_U24 ( .A(Midori_rounds_n1258), .Z(Midori_rounds_n1252)
         );
  BUF_X1 Midori_rounds_U23 ( .A(Midori_rounds_n2064), .Z(Midori_rounds_n1254)
         );
  INV_X1 Midori_rounds_U22 ( .A(Midori_rounds_n1275), .ZN(Midori_rounds_n1272)
         );
  INV_X1 Midori_rounds_U21 ( .A(Midori_rounds_n1275), .ZN(Midori_rounds_n1273)
         );
  INV_X1 Midori_rounds_U20 ( .A(Midori_rounds_n1275), .ZN(Midori_rounds_n1271)
         );
  BUF_X1 Midori_rounds_U19 ( .A(Midori_rounds_n1247), .Z(Midori_rounds_n1244)
         );
  INV_X1 Midori_rounds_U18 ( .A(Midori_rounds_n1275), .ZN(Midori_rounds_n1274)
         );
  INV_X1 Midori_rounds_U17 ( .A(Midori_rounds_n1275), .ZN(Midori_rounds_n1270)
         );
  BUF_X1 Midori_rounds_U16 ( .A(Midori_rounds_n1281), .Z(Midori_rounds_n1280)
         );
  BUF_X1 Midori_rounds_U15 ( .A(Midori_rounds_n1265), .Z(Midori_rounds_n1261)
         );
  BUF_X1 Midori_rounds_U14 ( .A(Midori_rounds_n1246), .Z(Midori_rounds_n1245)
         );
  BUF_X1 Midori_rounds_U13 ( .A(Midori_rounds_n1490), .Z(Midori_rounds_n1250)
         );
  BUF_X1 Midori_rounds_U12 ( .A(Midori_rounds_n1262), .Z(Midori_rounds_n1260)
         );
  BUF_X1 Midori_rounds_U11 ( .A(Midori_rounds_n1281), .Z(Midori_rounds_n1276)
         );
  INV_X1 Midori_rounds_U10 ( .A(Midori_rounds_n1276), .ZN(Midori_rounds_n1267)
         );
  BUF_X1 Midori_rounds_U9 ( .A(Midori_rounds_n1281), .Z(Midori_rounds_n1275)
         );
  BUF_X1 Midori_rounds_U8 ( .A(Midori_rounds_n1281), .Z(Midori_rounds_n1277)
         );
  BUF_X1 Midori_rounds_U7 ( .A(Midori_rounds_n1277), .Z(Midori_rounds_n1278)
         );
  OR2_X1 Midori_rounds_U6 ( .A1(enc_dec), .A2(reset), .ZN(Midori_rounds_n2066)
         );
  INV_X4 Midori_rounds_U5 ( .A(round_Signal[0]), .ZN(Midori_rounds_n1281) );
  XOR2_X1 Midori_rounds_U4 ( .A(Midori_rounds_n1241), .B(
        Midori_rounds_round_Constant[5]), .Z(Midori_rounds_n2048) );
  AOI22_X1 Midori_rounds_U3 ( .A1(round_Signal[0]), .A2(Key1[20]), .B1(
        Midori_rounds_n1277), .B2(Key1[84]), .ZN(Midori_rounds_n1241) );
  NAND3_X1 Midori_rounds_constant_MUX_U78 ( .A1(Midori_rounds_constant_MUX_n70), .A2(Midori_rounds_constant_MUX_n69), .A3(Midori_rounds_constant_MUX_n68), 
        .ZN(Midori_rounds_round_Constant[9]) );
  INV_X1 Midori_rounds_constant_MUX_U77 ( .A(Midori_rounds_constant_MUX_n67), 
        .ZN(Midori_rounds_constant_MUX_n70) );
  OR3_X1 Midori_rounds_constant_MUX_U76 ( .A1(Midori_rounds_constant_MUX_n66), 
        .A2(Midori_rounds_constant_MUX_n65), .A3(
        Midori_rounds_constant_MUX_n64), .ZN(Midori_rounds_round_Constant[8])
         );
  NAND4_X1 Midori_rounds_constant_MUX_U75 ( .A1(Midori_rounds_constant_MUX_n63), .A2(Midori_rounds_constant_MUX_n62), .A3(Midori_rounds_constant_MUX_n61), 
        .A4(Midori_rounds_constant_MUX_n60), .ZN(
        Midori_rounds_round_Constant[7]) );
  NAND3_X1 Midori_rounds_constant_MUX_U74 ( .A1(Midori_rounds_constant_MUX_n59), .A2(Midori_rounds_constant_MUX_n58), .A3(Midori_rounds_constant_MUX_n69), 
        .ZN(Midori_rounds_round_Constant[6]) );
  NAND2_X1 Midori_rounds_constant_MUX_U73 ( .A1(Midori_rounds_constant_MUX_n54), .A2(Midori_rounds_constant_MUX_n55), .ZN(Midori_rounds_round_Constant[4]) );
  NOR3_X1 Midori_rounds_constant_MUX_U72 ( .A1(Midori_rounds_constant_MUX_n53), 
        .A2(Midori_rounds_constant_MUX_n66), .A3(
        Midori_rounds_constant_MUX_n52), .ZN(Midori_rounds_constant_MUX_n55)
         );
  NAND2_X1 Midori_rounds_constant_MUX_U71 ( .A1(Midori_rounds_constant_MUX_n51), .A2(Midori_rounds_constant_MUX_n50), .ZN(Midori_rounds_round_Constant[3]) );
  NOR4_X1 Midori_rounds_constant_MUX_U70 ( .A1(Midori_rounds_constant_MUX_n49), 
        .A2(Midori_rounds_constant_MUX_n64), .A3(
        Midori_rounds_constant_MUX_n48), .A4(Midori_rounds_constant_MUX_n53), 
        .ZN(Midori_rounds_constant_MUX_n50) );
  NAND3_X1 Midori_rounds_constant_MUX_U69 ( .A1(Midori_rounds_constant_MUX_n61), .A2(Midori_rounds_constant_MUX_n47), .A3(Midori_rounds_constant_MUX_n69), 
        .ZN(Midori_rounds_round_Constant[2]) );
  NOR2_X1 Midori_rounds_constant_MUX_U68 ( .A1(Midori_rounds_constant_MUX_n64), 
        .A2(Midori_rounds_constant_MUX_n56), .ZN(
        Midori_rounds_constant_MUX_n69) );
  NAND4_X1 Midori_rounds_constant_MUX_U67 ( .A1(Midori_rounds_constant_MUX_n51), .A2(Midori_rounds_constant_MUX_n46), .A3(Midori_rounds_constant_MUX_n61), 
        .A4(Midori_rounds_constant_MUX_n45), .ZN(
        Midori_rounds_round_Constant[1]) );
  NOR3_X1 Midori_rounds_constant_MUX_U66 ( .A1(Midori_rounds_constant_MUX_n44), 
        .A2(Midori_rounds_constant_MUX_n48), .A3(
        Midori_rounds_constant_MUX_n56), .ZN(Midori_rounds_constant_MUX_n45)
         );
  OAI22_X1 Midori_rounds_constant_MUX_U65 ( .A1(Midori_rounds_constant_MUX_n43), .A2(Midori_rounds_constant_MUX_n42), .B1(Midori_rounds_constant_MUX_n41), 
        .B2(Midori_rounds_constant_MUX_n40), .ZN(
        Midori_rounds_constant_MUX_n56) );
  NAND3_X1 Midori_rounds_constant_MUX_U64 ( .A1(Midori_rounds_constant_MUX_n51), .A2(Midori_rounds_constant_MUX_n59), .A3(Midori_rounds_constant_MUX_n39), 
        .ZN(Midori_rounds_round_Constant[15]) );
  NAND3_X1 Midori_rounds_constant_MUX_U63 ( .A1(Midori_rounds_constant_MUX_n63), .A2(Midori_rounds_constant_MUX_n38), .A3(Midori_rounds_constant_MUX_n54), 
        .ZN(Midori_rounds_round_Constant[14]) );
  NOR2_X1 Midori_rounds_constant_MUX_U62 ( .A1(Midori_rounds_constant_MUX_n44), 
        .A2(Midori_rounds_constant_MUX_n65), .ZN(
        Midori_rounds_constant_MUX_n54) );
  INV_X1 Midori_rounds_constant_MUX_U61 ( .A(Midori_rounds_constant_MUX_n37), 
        .ZN(Midori_rounds_constant_MUX_n65) );
  INV_X1 Midori_rounds_constant_MUX_U60 ( .A(Midori_rounds_constant_MUX_n53), 
        .ZN(Midori_rounds_constant_MUX_n63) );
  OAI22_X1 Midori_rounds_constant_MUX_U59 ( .A1(Midori_rounds_constant_MUX_n36), .A2(Midori_rounds_constant_MUX_n35), .B1(Midori_rounds_constant_MUX_n34), 
        .B2(Midori_rounds_constant_MUX_n33), .ZN(
        Midori_rounds_constant_MUX_n53) );
  NAND4_X1 Midori_rounds_constant_MUX_U58 ( .A1(Midori_rounds_constant_MUX_n38), .A2(Midori_rounds_constant_MUX_n32), .A3(Midori_rounds_constant_MUX_n61), 
        .A4(Midori_rounds_constant_MUX_n31), .ZN(
        Midori_rounds_round_Constant[13]) );
  NOR2_X1 Midori_rounds_constant_MUX_U57 ( .A1(Midori_rounds_constant_MUX_n49), 
        .A2(Midori_rounds_constant_MUX_n30), .ZN(
        Midori_rounds_constant_MUX_n61) );
  AOI21_X1 Midori_rounds_constant_MUX_U56 ( .B1(Midori_rounds_constant_MUX_n29), .B2(Midori_rounds_constant_MUX_n28), .A(Midori_rounds_constant_MUX_n34), 
        .ZN(Midori_rounds_constant_MUX_n49) );
  INV_X1 Midori_rounds_constant_MUX_U55 ( .A(Midori_rounds_constant_MUX_n52), 
        .ZN(Midori_rounds_constant_MUX_n32) );
  INV_X1 Midori_rounds_constant_MUX_U54 ( .A(Midori_rounds_constant_MUX_n27), 
        .ZN(Midori_rounds_constant_MUX_n38) );
  NAND3_X1 Midori_rounds_constant_MUX_U53 ( .A1(Midori_rounds_constant_MUX_n37), .A2(Midori_rounds_constant_MUX_n62), .A3(Midori_rounds_constant_MUX_n58), 
        .ZN(Midori_rounds_round_Constant[12]) );
  NOR2_X1 Midori_rounds_constant_MUX_U52 ( .A1(Midori_rounds_constant_MUX_n27), 
        .A2(Midori_rounds_constant_MUX_n48), .ZN(
        Midori_rounds_constant_MUX_n58) );
  NOR3_X1 Midori_rounds_constant_MUX_U51 ( .A1(Midori_rounds_constant_MUX_n67), 
        .A2(Midori_rounds_constant_MUX_n57), .A3(
        Midori_rounds_constant_MUX_n30), .ZN(Midori_rounds_constant_MUX_n37)
         );
  OAI211_X1 Midori_rounds_constant_MUX_U50 ( .C1(
        Midori_rounds_constant_MUX_n33), .C2(Midori_rounds_constant_MUX_n41), 
        .A(Midori_rounds_constant_MUX_n26), .B(Midori_rounds_constant_MUX_n59), 
        .ZN(Midori_rounds_constant_MUX_n57) );
  INV_X1 Midori_rounds_constant_MUX_U49 ( .A(Midori_rounds_constant_MUX_n25), 
        .ZN(Midori_rounds_constant_MUX_n59) );
  OAI22_X1 Midori_rounds_constant_MUX_U48 ( .A1(Midori_rounds_constant_MUX_n36), .A2(Midori_rounds_constant_MUX_n24), .B1(Midori_rounds_constant_MUX_n34), 
        .B2(Midori_rounds_constant_MUX_n43), .ZN(
        Midori_rounds_constant_MUX_n25) );
  OR2_X1 Midori_rounds_constant_MUX_U47 ( .A1(Midori_rounds_constant_MUX_n42), 
        .A2(Midori_rounds_constant_MUX_n28), .ZN(
        Midori_rounds_constant_MUX_n26) );
  INV_X1 Midori_rounds_constant_MUX_U46 ( .A(Midori_rounds_constant_MUX_n60), 
        .ZN(Midori_rounds_round_Constant[11]) );
  NOR3_X1 Midori_rounds_constant_MUX_U45 ( .A1(Midori_rounds_constant_MUX_n67), 
        .A2(Midori_rounds_constant_MUX_n27), .A3(
        Midori_rounds_constant_MUX_n64), .ZN(Midori_rounds_constant_MUX_n60)
         );
  NOR3_X1 Midori_rounds_constant_MUX_U44 ( .A1(Midori_rounds_constant_MUX_n36), 
        .A2(Midori_rounds_constant_MUX_n23), .A3(round_Signal[3]), .ZN(
        Midori_rounds_constant_MUX_n64) );
  OAI211_X1 Midori_rounds_constant_MUX_U43 ( .C1(
        Midori_rounds_constant_MUX_n34), .C2(Midori_rounds_constant_MUX_n24), 
        .A(Midori_rounds_constant_MUX_n22), .B(Midori_rounds_constant_MUX_n51), 
        .ZN(Midori_rounds_constant_MUX_n27) );
  INV_X1 Midori_rounds_constant_MUX_U42 ( .A(Midori_rounds_constant_MUX_n21), 
        .ZN(Midori_rounds_constant_MUX_n51) );
  OAI22_X1 Midori_rounds_constant_MUX_U41 ( .A1(Midori_rounds_constant_MUX_n36), .A2(Midori_rounds_constant_MUX_n33), .B1(Midori_rounds_constant_MUX_n35), 
        .B2(Midori_rounds_constant_MUX_n34), .ZN(
        Midori_rounds_constant_MUX_n21) );
  OR2_X1 Midori_rounds_constant_MUX_U40 ( .A1(Midori_rounds_constant_MUX_n36), 
        .A2(Midori_rounds_constant_MUX_n43), .ZN(
        Midori_rounds_constant_MUX_n22) );
  NAND2_X1 Midori_rounds_constant_MUX_U39 ( .A1(round_Signal[2]), .A2(
        Midori_rounds_constant_MUX_n10), .ZN(Midori_rounds_constant_MUX_n36)
         );
  NAND2_X1 Midori_rounds_constant_MUX_U38 ( .A1(Midori_rounds_constant_MUX_n46), .A2(Midori_rounds_constant_MUX_n39), .ZN(Midori_rounds_round_Constant[10])
         );
  NOR3_X1 Midori_rounds_constant_MUX_U37 ( .A1(Midori_rounds_constant_MUX_n67), 
        .A2(Midori_rounds_constant_MUX_n52), .A3(
        Midori_rounds_constant_MUX_n20), .ZN(Midori_rounds_constant_MUX_n39)
         );
  OAI21_X1 Midori_rounds_constant_MUX_U36 ( .B1(Midori_rounds_constant_MUX_n35), .B2(Midori_rounds_constant_MUX_n42), .A(Midori_rounds_constant_MUX_n19), 
        .ZN(Midori_rounds_constant_MUX_n67) );
  OAI211_X1 Midori_rounds_constant_MUX_U35 ( .C1(
        Midori_rounds_constant_MUX_n18), .C2(Midori_rounds_constant_MUX_n10), 
        .A(round_Signal[2]), .B(Midori_rounds_constant_MUX_n17), .ZN(
        Midori_rounds_constant_MUX_n19) );
  INV_X1 Midori_rounds_constant_MUX_U34 ( .A(Midori_rounds_constant_MUX_n66), 
        .ZN(Midori_rounds_constant_MUX_n46) );
  NAND4_X1 Midori_rounds_constant_MUX_U33 ( .A1(Midori_rounds_constant_MUX_n16), .A2(Midori_rounds_constant_MUX_n62), .A3(Midori_rounds_constant_MUX_n47), 
        .A4(Midori_rounds_constant_MUX_n31), .ZN(
        Midori_rounds_round_Constant[0]) );
  INV_X1 Midori_rounds_constant_MUX_U32 ( .A(Midori_rounds_constant_MUX_n44), 
        .ZN(Midori_rounds_constant_MUX_n31) );
  AOI221_X1 Midori_rounds_constant_MUX_U31 ( .B1(round_Signal[3]), .B2(
        Midori_rounds_constant_MUX_n18), .C1(Midori_rounds_constant_MUX_n15), 
        .C2(enc_dec), .A(Midori_rounds_constant_MUX_n68), .ZN(
        Midori_rounds_constant_MUX_n44) );
  OR2_X1 Midori_rounds_constant_MUX_U30 ( .A1(Midori_rounds_constant_MUX_n23), 
        .A2(Midori_rounds_constant_MUX_n34), .ZN(
        Midori_rounds_constant_MUX_n68) );
  NAND2_X1 Midori_rounds_constant_MUX_U29 ( .A1(Midori_rounds_constant_MUX_n14), .A2(Midori_rounds_constant_MUX_n10), .ZN(Midori_rounds_constant_MUX_n34) );
  NOR2_X1 Midori_rounds_constant_MUX_U28 ( .A1(Midori_rounds_constant_MUX_n52), 
        .A2(Midori_rounds_constant_MUX_n48), .ZN(
        Midori_rounds_constant_MUX_n47) );
  OAI22_X1 Midori_rounds_constant_MUX_U27 ( .A1(Midori_rounds_constant_MUX_n24), .A2(Midori_rounds_constant_MUX_n41), .B1(Midori_rounds_constant_MUX_n42), 
        .B2(Midori_rounds_constant_MUX_n13), .ZN(
        Midori_rounds_constant_MUX_n48) );
  OAI22_X1 Midori_rounds_constant_MUX_U26 ( .A1(Midori_rounds_constant_MUX_n43), .A2(Midori_rounds_constant_MUX_n41), .B1(Midori_rounds_constant_MUX_n42), 
        .B2(Midori_rounds_constant_MUX_n40), .ZN(
        Midori_rounds_constant_MUX_n52) );
  NAND2_X1 Midori_rounds_constant_MUX_U25 ( .A1(round_Signal[1]), .A2(
        Midori_rounds_constant_MUX_n12), .ZN(Midori_rounds_constant_MUX_n40)
         );
  NOR2_X1 Midori_rounds_constant_MUX_U24 ( .A1(round_Signal[3]), .A2(enc_dec), 
        .ZN(Midori_rounds_constant_MUX_n12) );
  NAND3_X1 Midori_rounds_constant_MUX_U23 ( .A1(round_Signal[3]), .A2(enc_dec), 
        .A3(Midori_rounds_constant_MUX_n23), .ZN(
        Midori_rounds_constant_MUX_n43) );
  NOR2_X1 Midori_rounds_constant_MUX_U22 ( .A1(Midori_rounds_constant_MUX_n66), 
        .A2(Midori_rounds_constant_MUX_n20), .ZN(
        Midori_rounds_constant_MUX_n62) );
  OAI22_X1 Midori_rounds_constant_MUX_U21 ( .A1(Midori_rounds_constant_MUX_n33), .A2(Midori_rounds_constant_MUX_n42), .B1(Midori_rounds_constant_MUX_n28), 
        .B2(Midori_rounds_constant_MUX_n41), .ZN(
        Midori_rounds_constant_MUX_n20) );
  NAND3_X1 Midori_rounds_constant_MUX_U20 ( .A1(round_Signal[1]), .A2(enc_dec), 
        .A3(Midori_rounds_constant_MUX_n15), .ZN(
        Midori_rounds_constant_MUX_n28) );
  NAND3_X1 Midori_rounds_constant_MUX_U19 ( .A1(Midori_rounds_constant_MUX_n23), .A2(Midori_rounds_constant_MUX_n18), .A3(round_Signal[3]), .ZN(
        Midori_rounds_constant_MUX_n33) );
  OAI22_X1 Midori_rounds_constant_MUX_U18 ( .A1(Midori_rounds_constant_MUX_n24), .A2(Midori_rounds_constant_MUX_n42), .B1(Midori_rounds_constant_MUX_n41), 
        .B2(Midori_rounds_constant_MUX_n13), .ZN(
        Midori_rounds_constant_MUX_n66) );
  NAND2_X1 Midori_rounds_constant_MUX_U17 ( .A1(enc_dec), .A2(
        Midori_rounds_constant_MUX_n17), .ZN(Midori_rounds_constant_MUX_n13)
         );
  NAND3_X1 Midori_rounds_constant_MUX_U16 ( .A1(Midori_rounds_constant_MUX_n15), .A2(Midori_rounds_constant_MUX_n23), .A3(Midori_rounds_constant_MUX_n18), 
        .ZN(Midori_rounds_constant_MUX_n24) );
  INV_X1 Midori_rounds_constant_MUX_U15 ( .A(Midori_rounds_constant_MUX_n30), 
        .ZN(Midori_rounds_constant_MUX_n16) );
  OAI22_X1 Midori_rounds_constant_MUX_U14 ( .A1(Midori_rounds_constant_MUX_n35), .A2(Midori_rounds_constant_MUX_n41), .B1(Midori_rounds_constant_MUX_n29), 
        .B2(Midori_rounds_constant_MUX_n42), .ZN(
        Midori_rounds_constant_MUX_n30) );
  NAND2_X1 Midori_rounds_constant_MUX_U13 ( .A1(Midori_rounds_constant_MUX_n14), .A2(Midori_rounds_constant_MUX_n11), .ZN(Midori_rounds_constant_MUX_n42) );
  INV_X1 Midori_rounds_constant_MUX_U12 ( .A(round_Signal[2]), .ZN(
        Midori_rounds_constant_MUX_n14) );
  NAND2_X1 Midori_rounds_constant_MUX_U11 ( .A1(Midori_rounds_constant_MUX_n18), .A2(Midori_rounds_constant_MUX_n17), .ZN(Midori_rounds_constant_MUX_n29) );
  NOR2_X1 Midori_rounds_constant_MUX_U10 ( .A1(Midori_rounds_constant_MUX_n15), 
        .A2(Midori_rounds_constant_MUX_n23), .ZN(
        Midori_rounds_constant_MUX_n17) );
  INV_X1 Midori_rounds_constant_MUX_U9 ( .A(enc_dec), .ZN(
        Midori_rounds_constant_MUX_n18) );
  NAND2_X1 Midori_rounds_constant_MUX_U8 ( .A1(Midori_rounds_constant_MUX_n11), 
        .A2(round_Signal[2]), .ZN(Midori_rounds_constant_MUX_n41) );
  NAND3_X1 Midori_rounds_constant_MUX_U7 ( .A1(Midori_rounds_constant_MUX_n15), 
        .A2(Midori_rounds_constant_MUX_n23), .A3(enc_dec), .ZN(
        Midori_rounds_constant_MUX_n35) );
  INV_X1 Midori_rounds_constant_MUX_U6 ( .A(round_Signal[1]), .ZN(
        Midori_rounds_constant_MUX_n23) );
  INV_X1 Midori_rounds_constant_MUX_U5 ( .A(round_Signal[3]), .ZN(
        Midori_rounds_constant_MUX_n15) );
  INV_X1 Midori_rounds_constant_MUX_U4 ( .A(Midori_rounds_n1267), .ZN(
        Midori_rounds_constant_MUX_n11) );
  INV_X1 Midori_rounds_constant_MUX_U3 ( .A(Midori_rounds_constant_MUX_n11), 
        .ZN(Midori_rounds_constant_MUX_n10) );
  NAND2_X1 Midori_rounds_constant_MUX_U2 ( .A1(Midori_rounds_constant_MUX_n55), 
        .A2(Midori_rounds_constant_MUX_n9), .ZN(
        Midori_rounds_round_Constant[5]) );
  NOR2_X1 Midori_rounds_constant_MUX_U1 ( .A1(Midori_rounds_constant_MUX_n57), 
        .A2(Midori_rounds_constant_MUX_n56), .ZN(Midori_rounds_constant_MUX_n9) );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_InAff_out3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_S1_InAff_out3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_InAff_out3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_S1_InAff_out3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_InAff_out3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_S1_InAff_out3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_InAff_out3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_0_S1_InAff_out3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_S1_InAff_out2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_rs1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_S1_InAff_out2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_rs1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_S1_InAff_out2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_rs1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_0_S1_InAff_out2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_3_), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_S1_InAff_out1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_rs1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_S1_InAff_out1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_rs1[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_S1_InAff_out1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_rs1[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_0_S1_InAff_out1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_3_), .QN() );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_InputAffine_U3 ( .A(
        Midori_rounds_sub_Sub_0_S1_InAff_out3[1]), .B(Midori_rounds_n919), .Z(
        Midori_rounds_sub_Sub_0_S1_InAff_out3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_InputAffine_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_InAff_out2[1]), .B(Midori_rounds_n855), .Z(
        Midori_rounds_sub_Sub_0_S1_InAff_out2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_InputAffine_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_InAff_out1[1]), .B(Midori_rounds_n806), .Z(
        Midori_rounds_sub_Sub_0_S1_InAff_out1[3]) );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_rs1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_rs1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_0__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_rs2[0]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_0__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[0]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_0__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_rs1[1]), .C2(Midori_rounds_sub_Sub_0_rs1[2]), 
        .A(Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_0__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_0__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_rs1[1]), .A2(Midori_rounds_sub_Sub_0_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_0__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_0_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_U3 ( .A(r[0]), 
        .B(r[1]), .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_3_), .B2(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[1]), .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_1__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[2]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_0_rs1[1]), .C2(Midori_rounds_sub_Sub_0_rs1[2]), 
        .A(Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_0_rs1[1]), .A2(Midori_rounds_sub_Sub_0_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_rs2[1]), .B(Midori_rounds_sub_Sub_0_rs2[0]), 
        .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_U1 ( .A(r[2]), .B(
        r[1]), .Z(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_3__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_rs2[0]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_3__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[3]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_3__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_3__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_3__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_3__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_0_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_U3 ( .A(r[2]), 
        .B(r[3]), .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[3]), .B2(
        Midori_rounds_sub_Sub_0_rs1[4]), .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_0_rs1[5]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_4__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[5]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_rs2[1]), .B(Midori_rounds_sub_Sub_0_rs2[0]), 
        .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_U1 ( .A(r[4]), .B(
        r[3]), .Z(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_6__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_rs2[0]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_6__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[6]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_6__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_rs1[4]), .C2(Midori_rounds_sub_Sub_0_rs1[5]), 
        .A(Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_6__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_6__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_rs1[4]), .A2(Midori_rounds_sub_Sub_0_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_6__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[7]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_0_rs1[4]), .C2(Midori_rounds_sub_Sub_0_rs1[5]), 
        .A(Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_rs1[4]), .A2(Midori_rounds_sub_Sub_0_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_0_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_U1 ( .A(r[4]), 
        .B(r[5]), .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_7__CF_Inst_n9) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_n21), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_n20), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[8]) );
  OAI21_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_U5 ( .B1(
        Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_3_), .B2(
        Midori_rounds_sub_Sub_0_rs1[1]), .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_n19), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_n20) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_0_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_n19) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_n18), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_n17), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_n21) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_rs2[1]), .B(r[5]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_n17) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_rs2[0]), .B(r[0]), .Z(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_8__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_9__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_rs2[2]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_9__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[9]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_9__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_rs1[1]), .C2(Midori_rounds_sub_Sub_0_rs1[2]), 
        .A(Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_9__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_9__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_rs1[1]), .A2(Midori_rounds_sub_Sub_0_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_9__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_U3 ( .A(r[6]), 
        .B(r[7]), .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[2]), .B1(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_10__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[11]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_0_rs1[1]), .C2(Midori_rounds_sub_Sub_0_rs1[2]), 
        .A(Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_0_rs1[1]), .A2(Midori_rounds_sub_Sub_0_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_rs2[3]), .B(Midori_rounds_sub_Sub_0_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_U1 ( .A(r[8]), 
        .B(r[7]), .Z(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_rs2[2]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[12]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_12__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_12__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_12__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_U3 ( .A(r[8]), 
        .B(r[9]), .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_0_rs1[5]), .B1(Midori_rounds_sub_Sub_0_rs1[4]), 
        .B2(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_13__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[14]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_rs2[3]), .B(Midori_rounds_sub_Sub_0_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_U1 ( .A(r[10]), 
        .B(r[9]), .Z(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_15__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_rs2[2]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_15__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[15]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_15__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_rs1[4]), .C2(Midori_rounds_sub_Sub_0_rs1[5]), 
        .A(Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_15__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_15__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_rs1[4]), .A2(Midori_rounds_sub_Sub_0_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_15__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[16]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_0_rs1[4]), .C2(Midori_rounds_sub_Sub_0_rs1[5]), 
        .A(Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_rs1[4]), .A2(Midori_rounds_sub_Sub_0_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_0_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_U1 ( .A(r[10]), 
        .B(r[11]), .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_16__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_U4 ( .A(r[6]), 
        .B(Midori_rounds_sub_Sub_0_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_n16) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_U3 ( .A(r[11]), 
        .B(Midori_rounds_sub_Sub_0_rs2[3]), .Z(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_n17) );
  AOI22_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_0_rs1[2]), .B1(Midori_rounds_sub_Sub_0_rs1[1]), 
        .B2(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_17__CF_Inst_n15) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_18__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_rs2[4]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_18__CF_Inst_n3), .Z(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_rs1[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_18__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_U2 ( .A(r[13]), 
        .B(r[12]), .Z(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_rs2[5]), .B(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_19__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_0_rs1[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_U4 ( .A(r[13]), 
        .B(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_U2 ( .A(r[14]), 
        .B(Midori_rounds_sub_Sub_0_rs1[0]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_rs2[4]), .B(Midori_rounds_sub_Sub_0_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_20__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_21__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_21__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_0_rs2[4]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[21]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_21__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_rs1[4]), .A2(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_U2 ( .A(r[15]), 
        .B(r[14]), .Z(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_rs2[5]), .B(Midori_rounds_sub_Sub_0_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_22__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[23]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_U4 ( .A(r[15]), 
        .B(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_U2 ( .A(r[16]), 
        .B(Midori_rounds_sub_Sub_0_S1_InAff_out3_reg[0]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_rs2[4]), .B(Midori_rounds_sub_Sub_0_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_23__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_24__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_24__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_0_rs2[4]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[24]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_rs1[4]), .A2(
        Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_24__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[25]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_rs1[4]), .A2(
        Midori_rounds_sub_Sub_0_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_U2 ( .A(r[17]), 
        .B(r[16]), .Z(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_rs2[5]), .B(Midori_rounds_sub_Sub_0_rs1[3]), 
        .ZN(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_0_rs1[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_U4 ( .A(r[17]), 
        .B(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_U2 ( .A(r[12]), 
        .B(Midori_rounds_sub_Sub_0_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_rs2[4]), .B(Midori_rounds_sub_Sub_0_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_0_S1_F_inst_Inst_26__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_1__Compression2_n2), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_1__Compression2_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_0_S1_F_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_0_S1_F_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[49]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result1[49]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[49]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_0__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_0__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[0]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_0__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_U2 ( .A(r[31]), 
        .B(r[30]), .Z(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_0_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_1__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_U2 ( .A(1'b0), .B(
        r[32]), .Z(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_U1 ( .A(1'b0), 
        .B(r[31]), .ZN(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_3__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_3__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_U2 ( .A(r[33]), 
        .B(r[32]), .Z(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_0_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_4__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[5]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_U2 ( .A(1'b0), .B(
        r[34]), .Z(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_U1 ( .A(1'b0), 
        .B(r[33]), .ZN(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_6__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_6__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[6]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_6__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_7__CF_Inst_U4 ( .A(1'b0), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_7__CF_Inst_n9), .Z(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_7__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_7__CF_Inst_n8), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_7__CF_Inst_n7), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_7__CF_Inst_n9) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_7__CF_Inst_n7) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_7__CF_Inst_U1 ( .A(r[34]), 
        .B(r[35]), .Z(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_7__CF_Inst_n8) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_U4 ( .A(r[35]), 
        .B(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_U2 ( .A(r[30]), 
        .B(Midori_rounds_sub_Sub_0_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_U1 ( .A(1'b0), .B(
        1'b0), .Z(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_8__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_9__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_9__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[9]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[1]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_U1 ( .A(r[18]), 
        .B(r[19]), .Z(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_10__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[11]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_U4 ( .A(r[19]), 
        .B(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_U2 ( .A(r[20]), 
        .B(Midori_rounds_sub_Sub_0_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_12__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[1]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_U1 ( .A(r[20]), 
        .B(r[21]), .Z(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_13__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[14]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_U4 ( .A(r[21]), 
        .B(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_U2 ( .A(r[22]), 
        .B(Midori_rounds_sub_Sub_0_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_15__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_15__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[15]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_U2 ( .A(r[23]), 
        .B(r[22]), .Z(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_0_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_n13), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_n12), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_n12) );
  INV_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[1]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_U2 ( .A(r[23]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_n13)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_U1 ( .A(r[18]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_17__CF_Inst_n15)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_18__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_18__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[18]) );
  AOI21_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_18__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_18__CF_Inst_n6) );
  OAI21_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_18__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_U3 ( .A(r[24]), 
        .B(r[25]), .ZN(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[2]), .B1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[1]), .B2(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_19__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[20]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[1]), .C2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_U1 ( .A(r[26]), 
        .B(r[25]), .Z(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_20__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_21__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_21__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[21]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_21__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_21__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_U3 ( .A(r[26]), 
        .B(r[27]), .ZN(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[2]), .B1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[1]), .B2(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_22__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[23]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_U1 ( .A(r[28]), 
        .B(r[27]), .Z(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_23__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_24__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_24__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[24]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_24__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[25]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[3]), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_n9), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_U1 ( .A(r[28]), 
        .B(r[29]), .ZN(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_25__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Out[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_U4 ( .A(r[24]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_n16)
         );
  XOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_U3 ( .A(r[29]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_n17)
         );
  AOI22_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[2]), .B1(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[48]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[48]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[48]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[50]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[50]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[50]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[51]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[51]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[51]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_0_S1_G_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_0_S1_G_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_InAff_out3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_S2_InAff_out3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_InAff_out3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_S2_InAff_out3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_InAff_out3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_S2_InAff_out3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_InAff_out3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_0_S2_InAff_out3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_S2_InAff_out2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_rs2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_S2_InAff_out2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_rs2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_S2_InAff_out2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_rs2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_0_S2_InAff_out2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_3_), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_S2_InAff_out1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_rs2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_S2_InAff_out1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_rs2[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_S2_InAff_out1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_rs2[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_0_S2_InAff_out1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_3_), .QN() );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_InputAffine_U3 ( .A(
        Midori_rounds_sub_Sub_0_S2_InAff_out3[1]), .B(Midori_rounds_n923), .Z(
        Midori_rounds_sub_Sub_0_S2_InAff_out3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_InputAffine_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_InAff_out2[1]), .B(Midori_rounds_n859), .Z(
        Midori_rounds_sub_Sub_0_S2_InAff_out2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_InputAffine_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_InAff_out1[1]), .B(Midori_rounds_n809), .Z(
        Midori_rounds_sub_Sub_0_S2_InAff_out1[3]) );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_rs2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_rs2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_0__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_rs1[0]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_0__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[0]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_0__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_rs2[1]), .C2(Midori_rounds_sub_Sub_0_rs2[2]), 
        .A(Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_0__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_0__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_rs2[1]), .A2(Midori_rounds_sub_Sub_0_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_0__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_0_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_U3 ( .A(r[36]), 
        .B(r[37]), .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_3_), .B2(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[1]), .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_1__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[2]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_0_rs2[1]), .C2(Midori_rounds_sub_Sub_0_rs2[2]), 
        .A(Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_0_rs2[1]), .A2(Midori_rounds_sub_Sub_0_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_rs1[1]), .B(Midori_rounds_sub_Sub_0_rs1[0]), 
        .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_U1 ( .A(r[38]), 
        .B(r[37]), .Z(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_3__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_rs1[0]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_3__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[3]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_3__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_3__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_3__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_3__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_0_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_U3 ( .A(r[38]), 
        .B(r[39]), .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[3]), .B2(
        Midori_rounds_sub_Sub_0_rs2[4]), .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_0_rs2[5]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_4__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[5]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_rs1[1]), .B(Midori_rounds_sub_Sub_0_rs1[0]), 
        .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_U1 ( .A(r[40]), 
        .B(r[39]), .Z(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_6__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_rs1[0]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_6__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[6]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_6__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_rs2[4]), .C2(Midori_rounds_sub_Sub_0_rs2[5]), 
        .A(Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_6__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_6__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_rs2[4]), .A2(Midori_rounds_sub_Sub_0_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_6__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[7]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_0_rs2[4]), .C2(Midori_rounds_sub_Sub_0_rs2[5]), 
        .A(Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_rs2[4]), .A2(Midori_rounds_sub_Sub_0_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_0_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_U1 ( .A(r[40]), 
        .B(r[41]), .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_7__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_n21), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_n20), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[8]) );
  OAI21_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_U5 ( .B1(
        Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_3_), .B2(
        Midori_rounds_sub_Sub_0_rs2[1]), .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_n19), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_n20) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_0_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_n19) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_n18), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_n17), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_n21) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_rs1[1]), .B(r[41]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_n17) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_rs1[0]), .B(r[36]), .Z(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_8__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_9__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_rs1[2]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_9__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[9]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_9__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_rs2[1]), .C2(Midori_rounds_sub_Sub_0_rs2[2]), 
        .A(Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_9__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_9__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_rs2[1]), .A2(Midori_rounds_sub_Sub_0_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_9__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_U3 ( .A(r[42]), 
        .B(r[43]), .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[2]), .B1(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[1]), .B2(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_10__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[11]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_0_rs2[1]), .C2(Midori_rounds_sub_Sub_0_rs2[2]), 
        .A(Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_0_rs2[1]), .A2(Midori_rounds_sub_Sub_0_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_rs1[3]), .B(Midori_rounds_sub_Sub_0_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_U1 ( .A(r[44]), 
        .B(r[43]), .Z(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_rs1[2]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[12]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_12__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_12__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_12__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_U3 ( .A(r[44]), 
        .B(r[45]), .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_0_rs2[5]), .B1(Midori_rounds_sub_Sub_0_rs2[4]), 
        .B2(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_13__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[14]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_rs1[3]), .B(Midori_rounds_sub_Sub_0_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_U1 ( .A(r[46]), 
        .B(r[45]), .Z(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_15__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_rs1[2]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_15__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[15]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_15__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_rs2[4]), .C2(Midori_rounds_sub_Sub_0_rs2[5]), 
        .A(Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_15__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_15__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_rs2[4]), .A2(Midori_rounds_sub_Sub_0_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_15__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[16]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_0_rs2[4]), .C2(Midori_rounds_sub_Sub_0_rs2[5]), 
        .A(Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_rs2[4]), .A2(Midori_rounds_sub_Sub_0_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_0_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_U1 ( .A(r[46]), 
        .B(r[47]), .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_16__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_U4 ( .A(r[42]), 
        .B(Midori_rounds_sub_Sub_0_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_n16) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_U3 ( .A(r[47]), 
        .B(Midori_rounds_sub_Sub_0_rs1[3]), .Z(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_n17) );
  AOI22_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_0_rs2[2]), .B1(Midori_rounds_sub_Sub_0_rs2[1]), 
        .B2(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_17__CF_Inst_n15) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_18__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_rs1[4]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_18__CF_Inst_n3), .Z(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_rs2[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_18__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_U2 ( .A(r[49]), 
        .B(r[48]), .Z(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_rs1[5]), .B(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_19__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_0_rs2[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_U4 ( .A(r[49]), 
        .B(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_U2 ( .A(r[50]), 
        .B(Midori_rounds_sub_Sub_0_rs2[0]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_rs1[4]), .B(Midori_rounds_sub_Sub_0_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_20__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_21__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_21__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_0_rs1[4]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[21]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_21__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_rs2[4]), .A2(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_U2 ( .A(r[51]), 
        .B(r[50]), .Z(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_rs1[5]), .B(Midori_rounds_sub_Sub_0_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_22__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[23]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_U4 ( .A(r[51]), 
        .B(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_U2 ( .A(r[52]), 
        .B(Midori_rounds_sub_Sub_0_S2_InAff_out3_reg[0]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_rs1[4]), .B(Midori_rounds_sub_Sub_0_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_23__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_24__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_24__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_0_rs1[4]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[24]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_rs2[4]), .A2(
        Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_24__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[25]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_rs2[4]), .A2(
        Midori_rounds_sub_Sub_0_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_U2 ( .A(r[53]), 
        .B(r[52]), .Z(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_rs1[5]), .B(Midori_rounds_sub_Sub_0_rs2[3]), 
        .ZN(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_0_rs2[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_U4 ( .A(r[53]), 
        .B(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_U2 ( .A(r[48]), 
        .B(Midori_rounds_sub_Sub_0_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_rs1[4]), .B(Midori_rounds_sub_Sub_0_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_0_S2_F_inst_Inst_26__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_1__Compression2_n2), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_1__Compression2_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_0_S2_F_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_0_S2_F_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[45]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result1[45]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[45]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_0__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_0__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[0]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_0__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_U2 ( .A(r[67]), 
        .B(r[66]), .Z(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_0_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_1__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_U2 ( .A(1'b0), .B(
        r[68]), .Z(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_U1 ( .A(1'b0), 
        .B(r[67]), .ZN(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_3__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_3__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_U2 ( .A(r[69]), 
        .B(r[68]), .Z(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_0_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_4__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[5]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_U2 ( .A(1'b0), .B(
        r[70]), .Z(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_U1 ( .A(1'b0), 
        .B(r[69]), .ZN(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_6__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_6__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[6]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_6__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_7__CF_Inst_U4 ( .A(1'b0), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_7__CF_Inst_n9), .Z(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_7__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_7__CF_Inst_n8), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_7__CF_Inst_n7), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_7__CF_Inst_n9) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_7__CF_Inst_n7) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_7__CF_Inst_U1 ( .A(r[70]), 
        .B(r[71]), .Z(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_7__CF_Inst_n8) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_U4 ( .A(r[71]), 
        .B(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_U2 ( .A(r[66]), 
        .B(Midori_rounds_sub_Sub_0_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_U1 ( .A(1'b0), .B(
        1'b0), .Z(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_8__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_9__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_9__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[9]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[1]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_U1 ( .A(r[54]), 
        .B(r[55]), .Z(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_10__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[11]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_U4 ( .A(r[55]), 
        .B(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_U2 ( .A(r[56]), 
        .B(Midori_rounds_sub_Sub_0_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_12__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[1]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_U1 ( .A(r[56]), 
        .B(r[57]), .Z(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_13__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[14]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_U4 ( .A(r[57]), 
        .B(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_U2 ( .A(r[58]), 
        .B(Midori_rounds_sub_Sub_0_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_15__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_15__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[15]) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_U2 ( .A(r[59]), 
        .B(r[58]), .Z(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_0_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_n13), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_n12), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_n12) );
  INV_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[1]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_U2 ( .A(r[59]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_n13)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_U1 ( .A(r[54]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_17__CF_Inst_n15)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_18__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_18__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[18]) );
  AOI21_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_18__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_18__CF_Inst_n6) );
  OAI21_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_18__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_U3 ( .A(r[60]), 
        .B(r[61]), .ZN(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[2]), .B1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[1]), .B2(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_19__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[20]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[1]), .C2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_U1 ( .A(r[62]), 
        .B(r[61]), .Z(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_20__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_21__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_21__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[21]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_21__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_21__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_U3 ( .A(r[62]), 
        .B(r[63]), .ZN(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[2]), .B1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[1]), .B2(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_22__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[23]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_U1 ( .A(r[64]), 
        .B(r[63]), .Z(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_23__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_24__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_24__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[24]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_24__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[25]) );
  OAI211_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[3]), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_n9), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_U1 ( .A(r[64]), 
        .B(r[65]), .ZN(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_25__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Out[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_U4 ( .A(r[60]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_n16)
         );
  XOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_U3 ( .A(r[65]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_n17)
         );
  AOI22_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[2]), .B1(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[44]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[44]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[44]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[46]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[46]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[46]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[47]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[47]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[47]) );
  XNOR2_X1 Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_0_S2_G_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_0_S2_G_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_InAff_out3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_S1_InAff_out3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_InAff_out3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_S1_InAff_out3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_InAff_out3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_S1_InAff_out3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_InAff_out3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_1_S1_InAff_out3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_S1_InAff_out2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_rs1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_S1_InAff_out2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_rs1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_S1_InAff_out2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_rs1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_1_S1_InAff_out2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_3_), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_S1_InAff_out1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_rs1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_S1_InAff_out1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_rs1[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_S1_InAff_out1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_rs1[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_1_S1_InAff_out1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_3_), .QN() );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_InputAffine_U3 ( .A(
        Midori_rounds_sub_Sub_1_S1_InAff_out3[1]), .B(Midori_rounds_n927), .Z(
        Midori_rounds_sub_Sub_1_S1_InAff_out3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_InputAffine_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_InAff_out2[1]), .B(Midori_rounds_n863), .Z(
        Midori_rounds_sub_Sub_1_S1_InAff_out2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_InputAffine_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_InAff_out1[1]), .B(Midori_rounds_n812), .Z(
        Midori_rounds_sub_Sub_1_S1_InAff_out1[3]) );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_rs1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_rs1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_0__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_rs2[0]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_0__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[0]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_0__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_rs1[1]), .C2(Midori_rounds_sub_Sub_1_rs1[2]), 
        .A(Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_0__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_0__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_rs1[1]), .A2(Midori_rounds_sub_Sub_1_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_0__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_1_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_U3 ( .A(r[0]), 
        .B(r[1]), .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_3_), .B2(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[1]), .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_1__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[2]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_1_rs1[1]), .C2(Midori_rounds_sub_Sub_1_rs1[2]), 
        .A(Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_1_rs1[1]), .A2(Midori_rounds_sub_Sub_1_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_rs2[1]), .B(Midori_rounds_sub_Sub_1_rs2[0]), 
        .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_U1 ( .A(r[2]), .B(
        r[1]), .Z(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_3__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_rs2[0]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_3__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[3]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_3__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_3__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_3__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_3__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_1_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_U3 ( .A(r[2]), 
        .B(r[3]), .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[3]), .B2(
        Midori_rounds_sub_Sub_1_rs1[4]), .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_1_rs1[5]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_4__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[5]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_rs2[1]), .B(Midori_rounds_sub_Sub_1_rs2[0]), 
        .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_U1 ( .A(r[4]), .B(
        r[3]), .Z(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_6__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_rs2[0]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_6__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[6]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_6__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_rs1[4]), .C2(Midori_rounds_sub_Sub_1_rs1[5]), 
        .A(Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_6__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_6__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_rs1[4]), .A2(Midori_rounds_sub_Sub_1_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_6__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[7]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_1_rs1[4]), .C2(Midori_rounds_sub_Sub_1_rs1[5]), 
        .A(Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_rs1[4]), .A2(Midori_rounds_sub_Sub_1_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_1_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_U1 ( .A(r[4]), 
        .B(r[5]), .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_7__CF_Inst_n9) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_n21), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_n20), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[8]) );
  OAI21_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_U5 ( .B1(
        Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_3_), .B2(
        Midori_rounds_sub_Sub_1_rs1[1]), .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_n19), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_n20) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_1_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_n19) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_n18), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_n17), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_n21) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_rs2[1]), .B(r[5]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_n17) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_rs2[0]), .B(r[0]), .Z(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_8__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_9__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_rs2[2]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_9__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[9]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_9__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_rs1[1]), .C2(Midori_rounds_sub_Sub_1_rs1[2]), 
        .A(Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_9__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_9__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_rs1[1]), .A2(Midori_rounds_sub_Sub_1_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_9__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_U3 ( .A(r[6]), 
        .B(r[7]), .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[2]), .B1(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_10__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[11]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_1_rs1[1]), .C2(Midori_rounds_sub_Sub_1_rs1[2]), 
        .A(Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_1_rs1[1]), .A2(Midori_rounds_sub_Sub_1_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_rs2[3]), .B(Midori_rounds_sub_Sub_1_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_U1 ( .A(r[8]), 
        .B(r[7]), .Z(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_rs2[2]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[12]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_12__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_12__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_12__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_U3 ( .A(r[8]), 
        .B(r[9]), .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_1_rs1[5]), .B1(Midori_rounds_sub_Sub_1_rs1[4]), 
        .B2(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_13__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[14]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_rs2[3]), .B(Midori_rounds_sub_Sub_1_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_U1 ( .A(r[10]), 
        .B(r[9]), .Z(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_15__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_rs2[2]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_15__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[15]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_15__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_rs1[4]), .C2(Midori_rounds_sub_Sub_1_rs1[5]), 
        .A(Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_15__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_15__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_rs1[4]), .A2(Midori_rounds_sub_Sub_1_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_15__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[16]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_1_rs1[4]), .C2(Midori_rounds_sub_Sub_1_rs1[5]), 
        .A(Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_rs1[4]), .A2(Midori_rounds_sub_Sub_1_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_1_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_U1 ( .A(r[10]), 
        .B(r[11]), .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_16__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_U4 ( .A(r[6]), 
        .B(Midori_rounds_sub_Sub_1_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_n16) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_U3 ( .A(r[11]), 
        .B(Midori_rounds_sub_Sub_1_rs2[3]), .Z(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_n17) );
  AOI22_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_1_rs1[2]), .B1(Midori_rounds_sub_Sub_1_rs1[1]), 
        .B2(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_17__CF_Inst_n15) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_18__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_rs2[4]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_18__CF_Inst_n3), .Z(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_rs1[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_18__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_U2 ( .A(r[13]), 
        .B(r[12]), .Z(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_rs2[5]), .B(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_19__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_1_rs1[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_U4 ( .A(r[13]), 
        .B(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_U2 ( .A(r[14]), 
        .B(Midori_rounds_sub_Sub_1_rs1[0]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_rs2[4]), .B(Midori_rounds_sub_Sub_1_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_20__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_21__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_21__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_1_rs2[4]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[21]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_21__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_rs1[4]), .A2(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_U2 ( .A(r[15]), 
        .B(r[14]), .Z(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_rs2[5]), .B(Midori_rounds_sub_Sub_1_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_22__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[23]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_U4 ( .A(r[15]), 
        .B(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_U2 ( .A(r[16]), 
        .B(Midori_rounds_sub_Sub_1_S1_InAff_out3_reg[0]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_rs2[4]), .B(Midori_rounds_sub_Sub_1_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_23__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_24__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_24__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_1_rs2[4]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[24]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_rs1[4]), .A2(
        Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_24__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[25]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_rs1[4]), .A2(
        Midori_rounds_sub_Sub_1_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_U2 ( .A(r[17]), 
        .B(r[16]), .Z(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_rs2[5]), .B(Midori_rounds_sub_Sub_1_rs1[3]), 
        .ZN(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_1_rs1[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_U4 ( .A(r[17]), 
        .B(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_U2 ( .A(r[12]), 
        .B(Midori_rounds_sub_Sub_1_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_rs2[4]), .B(Midori_rounds_sub_Sub_1_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_1_S1_F_inst_Inst_26__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_1__Compression2_n2), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_1__Compression2_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_1_S1_F_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_1_S1_F_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result1[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_0__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_0__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[0]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_0__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_U2 ( .A(r[31]), 
        .B(r[30]), .Z(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_1_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_1__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_U2 ( .A(1'b0), .B(
        r[32]), .Z(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_U1 ( .A(1'b0), 
        .B(r[31]), .ZN(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_3__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_3__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_U2 ( .A(r[33]), 
        .B(r[32]), .Z(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_1_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_4__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[5]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_U2 ( .A(1'b0), .B(
        r[34]), .Z(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_U1 ( .A(1'b0), 
        .B(r[33]), .ZN(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_6__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_6__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[6]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_6__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_7__CF_Inst_U4 ( .A(1'b0), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_7__CF_Inst_n9), .Z(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_7__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_7__CF_Inst_n8), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_7__CF_Inst_n7), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_7__CF_Inst_n9) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_7__CF_Inst_n7) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_7__CF_Inst_U1 ( .A(r[34]), 
        .B(r[35]), .Z(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_7__CF_Inst_n8) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_U4 ( .A(r[35]), 
        .B(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_U2 ( .A(r[30]), 
        .B(Midori_rounds_sub_Sub_1_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_U1 ( .A(1'b0), .B(
        1'b0), .Z(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_8__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_9__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_9__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[9]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[1]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_U1 ( .A(r[18]), 
        .B(r[19]), .Z(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_10__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[11]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_U4 ( .A(r[19]), 
        .B(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_U2 ( .A(r[20]), 
        .B(Midori_rounds_sub_Sub_1_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_12__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[1]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_U1 ( .A(r[20]), 
        .B(r[21]), .Z(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_13__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[14]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_U4 ( .A(r[21]), 
        .B(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_U2 ( .A(r[22]), 
        .B(Midori_rounds_sub_Sub_1_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_15__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_15__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[15]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_U2 ( .A(r[23]), 
        .B(r[22]), .Z(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_1_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_n13), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_n12), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_n12) );
  INV_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[1]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_U2 ( .A(r[23]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_n13)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_U1 ( .A(r[18]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_17__CF_Inst_n15)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_18__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_18__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[18]) );
  AOI21_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_18__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_18__CF_Inst_n6) );
  OAI21_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_18__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_U3 ( .A(r[24]), 
        .B(r[25]), .ZN(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[2]), .B1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[1]), .B2(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_19__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[20]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[1]), .C2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_U1 ( .A(r[26]), 
        .B(r[25]), .Z(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_20__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_21__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_21__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[21]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_21__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_21__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_U3 ( .A(r[26]), 
        .B(r[27]), .ZN(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[2]), .B1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[1]), .B2(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_22__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[23]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_U1 ( .A(r[28]), 
        .B(r[27]), .Z(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_23__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_24__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_24__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[24]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_24__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[25]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[3]), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_n9), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_U1 ( .A(r[28]), 
        .B(r[29]), .ZN(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_25__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Out[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_U4 ( .A(r[24]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_n16)
         );
  XOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_U3 ( .A(r[29]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_n17)
         );
  AOI22_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[2]), .B1(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[8]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[8]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[8]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[11]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_1_S1_G_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_1_S1_G_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_InAff_out3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_S2_InAff_out3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_InAff_out3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_S2_InAff_out3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_InAff_out3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_S2_InAff_out3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_InAff_out3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_1_S2_InAff_out3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_S2_InAff_out2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_rs2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_S2_InAff_out2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_rs2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_S2_InAff_out2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_rs2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_1_S2_InAff_out2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_3_), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_S2_InAff_out1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_rs2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_S2_InAff_out1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_rs2[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_S2_InAff_out1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_rs2[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_1_S2_InAff_out1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_3_), .QN() );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_InputAffine_U3 ( .A(
        Midori_rounds_sub_Sub_1_S2_InAff_out3[1]), .B(Midori_rounds_n931), .Z(
        Midori_rounds_sub_Sub_1_S2_InAff_out3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_InputAffine_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_InAff_out2[1]), .B(Midori_rounds_n867), .Z(
        Midori_rounds_sub_Sub_1_S2_InAff_out2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_InputAffine_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_InAff_out1[1]), .B(Midori_rounds_n815), .Z(
        Midori_rounds_sub_Sub_1_S2_InAff_out1[3]) );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_rs2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_rs2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_0__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_rs1[0]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_0__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[0]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_0__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_rs2[1]), .C2(Midori_rounds_sub_Sub_1_rs2[2]), 
        .A(Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_0__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_0__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_rs2[1]), .A2(Midori_rounds_sub_Sub_1_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_0__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_1_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_U3 ( .A(r[36]), 
        .B(r[37]), .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_3_), .B2(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[1]), .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_1__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[2]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_1_rs2[1]), .C2(Midori_rounds_sub_Sub_1_rs2[2]), 
        .A(Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_1_rs2[1]), .A2(Midori_rounds_sub_Sub_1_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_rs1[1]), .B(Midori_rounds_sub_Sub_1_rs1[0]), 
        .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_U1 ( .A(r[38]), 
        .B(r[37]), .Z(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_3__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_rs1[0]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_3__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[3]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_3__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_3__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_3__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_3__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_1_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_U3 ( .A(r[38]), 
        .B(r[39]), .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[3]), .B2(
        Midori_rounds_sub_Sub_1_rs2[4]), .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_1_rs2[5]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_4__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[5]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_rs1[1]), .B(Midori_rounds_sub_Sub_1_rs1[0]), 
        .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_U1 ( .A(r[40]), 
        .B(r[39]), .Z(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_6__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_rs1[0]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_6__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[6]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_6__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_rs2[4]), .C2(Midori_rounds_sub_Sub_1_rs2[5]), 
        .A(Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_6__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_6__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_rs2[4]), .A2(Midori_rounds_sub_Sub_1_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_6__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[7]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_1_rs2[4]), .C2(Midori_rounds_sub_Sub_1_rs2[5]), 
        .A(Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_rs2[4]), .A2(Midori_rounds_sub_Sub_1_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_1_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_U1 ( .A(r[40]), 
        .B(r[41]), .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_7__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_n21), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_n20), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[8]) );
  OAI21_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_U5 ( .B1(
        Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_3_), .B2(
        Midori_rounds_sub_Sub_1_rs2[1]), .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_n19), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_n20) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_1_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_n19) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_n18), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_n17), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_n21) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_rs1[1]), .B(r[41]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_n17) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_rs1[0]), .B(r[36]), .Z(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_8__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_9__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_rs1[2]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_9__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[9]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_9__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_rs2[1]), .C2(Midori_rounds_sub_Sub_1_rs2[2]), 
        .A(Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_9__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_9__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_rs2[1]), .A2(Midori_rounds_sub_Sub_1_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_9__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_U3 ( .A(r[42]), 
        .B(r[43]), .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[2]), .B1(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[1]), .B2(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_10__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[11]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_1_rs2[1]), .C2(Midori_rounds_sub_Sub_1_rs2[2]), 
        .A(Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_1_rs2[1]), .A2(Midori_rounds_sub_Sub_1_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_rs1[3]), .B(Midori_rounds_sub_Sub_1_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_U1 ( .A(r[44]), 
        .B(r[43]), .Z(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_rs1[2]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[12]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_12__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_12__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_12__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_U3 ( .A(r[44]), 
        .B(r[45]), .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_1_rs2[5]), .B1(Midori_rounds_sub_Sub_1_rs2[4]), 
        .B2(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_13__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[14]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_rs1[3]), .B(Midori_rounds_sub_Sub_1_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_U1 ( .A(r[46]), 
        .B(r[45]), .Z(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_15__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_rs1[2]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_15__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[15]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_15__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_rs2[4]), .C2(Midori_rounds_sub_Sub_1_rs2[5]), 
        .A(Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_15__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_15__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_rs2[4]), .A2(Midori_rounds_sub_Sub_1_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_15__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[16]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_1_rs2[4]), .C2(Midori_rounds_sub_Sub_1_rs2[5]), 
        .A(Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_rs2[4]), .A2(Midori_rounds_sub_Sub_1_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_1_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_U1 ( .A(r[46]), 
        .B(r[47]), .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_16__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_U4 ( .A(r[42]), 
        .B(Midori_rounds_sub_Sub_1_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_n16) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_U3 ( .A(r[47]), 
        .B(Midori_rounds_sub_Sub_1_rs1[3]), .Z(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_n17) );
  AOI22_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_1_rs2[2]), .B1(Midori_rounds_sub_Sub_1_rs2[1]), 
        .B2(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_17__CF_Inst_n15) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_18__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_rs1[4]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_18__CF_Inst_n3), .Z(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_rs2[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_18__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_U2 ( .A(r[49]), 
        .B(r[48]), .Z(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_rs1[5]), .B(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_19__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_1_rs2[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_U4 ( .A(r[49]), 
        .B(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_U2 ( .A(r[50]), 
        .B(Midori_rounds_sub_Sub_1_rs2[0]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_rs1[4]), .B(Midori_rounds_sub_Sub_1_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_20__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_21__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_21__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_1_rs1[4]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[21]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_21__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_rs2[4]), .A2(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_U2 ( .A(r[51]), 
        .B(r[50]), .Z(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_rs1[5]), .B(Midori_rounds_sub_Sub_1_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_22__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[23]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_U4 ( .A(r[51]), 
        .B(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_U2 ( .A(r[52]), 
        .B(Midori_rounds_sub_Sub_1_S2_InAff_out3_reg[0]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_rs1[4]), .B(Midori_rounds_sub_Sub_1_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_23__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_24__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_24__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_1_rs1[4]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[24]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_rs2[4]), .A2(
        Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_24__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[25]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_rs2[4]), .A2(
        Midori_rounds_sub_Sub_1_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_U2 ( .A(r[53]), 
        .B(r[52]), .Z(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_rs1[5]), .B(Midori_rounds_sub_Sub_1_rs2[3]), 
        .ZN(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_1_rs2[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_U4 ( .A(r[53]), 
        .B(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_U2 ( .A(r[48]), 
        .B(Midori_rounds_sub_Sub_1_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_rs1[4]), .B(Midori_rounds_sub_Sub_1_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_1_S2_F_inst_Inst_26__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_1__Compression2_n2), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_1__Compression2_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_1_S2_F_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_1_S2_F_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result1[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_0__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_0__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[0]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_0__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_U2 ( .A(r[67]), 
        .B(r[66]), .Z(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_1_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_1__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_U2 ( .A(1'b0), .B(
        r[68]), .Z(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_U1 ( .A(1'b0), 
        .B(r[67]), .ZN(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_3__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_3__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_U2 ( .A(r[69]), 
        .B(r[68]), .Z(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_1_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_4__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[5]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_U2 ( .A(1'b0), .B(
        r[70]), .Z(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_U1 ( .A(1'b0), 
        .B(r[69]), .ZN(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_6__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_6__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[6]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_6__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_7__CF_Inst_U4 ( .A(1'b0), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_7__CF_Inst_n9), .Z(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_7__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_7__CF_Inst_n8), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_7__CF_Inst_n7), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_7__CF_Inst_n9) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_7__CF_Inst_n7) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_7__CF_Inst_U1 ( .A(r[70]), 
        .B(r[71]), .Z(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_7__CF_Inst_n8) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_U4 ( .A(r[71]), 
        .B(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_U2 ( .A(r[66]), 
        .B(Midori_rounds_sub_Sub_1_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_U1 ( .A(1'b0), .B(
        1'b0), .Z(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_8__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_9__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_9__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[9]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[1]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_U1 ( .A(r[54]), 
        .B(r[55]), .Z(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_10__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[11]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_U4 ( .A(r[55]), 
        .B(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_U2 ( .A(r[56]), 
        .B(Midori_rounds_sub_Sub_1_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_12__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[1]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_U1 ( .A(r[56]), 
        .B(r[57]), .Z(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_13__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[14]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_U4 ( .A(r[57]), 
        .B(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_U2 ( .A(r[58]), 
        .B(Midori_rounds_sub_Sub_1_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_15__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_15__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[15]) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_U2 ( .A(r[59]), 
        .B(r[58]), .Z(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_1_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_n13), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_n12), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_n12) );
  INV_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[1]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_U2 ( .A(r[59]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_n13)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_U1 ( .A(r[54]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_17__CF_Inst_n15)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_18__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_18__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[18]) );
  AOI21_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_18__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_18__CF_Inst_n6) );
  OAI21_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_18__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_U3 ( .A(r[60]), 
        .B(r[61]), .ZN(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[2]), .B1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[1]), .B2(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_19__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[20]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[1]), .C2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_U1 ( .A(r[62]), 
        .B(r[61]), .Z(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_20__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_21__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_21__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[21]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_21__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_21__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_U3 ( .A(r[62]), 
        .B(r[63]), .ZN(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[2]), .B1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[1]), .B2(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_22__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[23]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_U1 ( .A(r[64]), 
        .B(r[63]), .Z(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_23__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_24__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_24__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[24]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_24__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[25]) );
  OAI211_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[3]), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_n9), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_U1 ( .A(r[64]), 
        .B(r[65]), .ZN(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_25__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Out[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_U4 ( .A(r[60]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_n16)
         );
  XOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_U3 ( .A(r[65]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_n17)
         );
  AOI22_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[2]), .B1(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[20]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[20]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[20]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[23]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[23]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[23]) );
  XNOR2_X1 Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_1_S2_G_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_1_S2_G_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_InAff_out3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_S1_InAff_out3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_InAff_out3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_S1_InAff_out3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_InAff_out3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_S1_InAff_out3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_InAff_out3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_2_S1_InAff_out3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_S1_InAff_out2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_rs1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_S1_InAff_out2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_rs1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_S1_InAff_out2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_rs1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_2_S1_InAff_out2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_3_), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_S1_InAff_out1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_rs1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_S1_InAff_out1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_rs1[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_S1_InAff_out1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_rs1[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_2_S1_InAff_out1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_3_), .QN() );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_InputAffine_U3 ( .A(
        Midori_rounds_sub_Sub_2_S1_InAff_out3[1]), .B(Midori_rounds_n935), .Z(
        Midori_rounds_sub_Sub_2_S1_InAff_out3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_InputAffine_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_InAff_out2[1]), .B(Midori_rounds_n871), .Z(
        Midori_rounds_sub_Sub_2_S1_InAff_out2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_InputAffine_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_InAff_out1[1]), .B(Midori_rounds_n818), .Z(
        Midori_rounds_sub_Sub_2_S1_InAff_out1[3]) );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_rs1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_rs1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_0__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_rs2[0]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_0__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[0]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_0__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_rs1[1]), .C2(Midori_rounds_sub_Sub_2_rs1[2]), 
        .A(Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_0__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_0__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_rs1[1]), .A2(Midori_rounds_sub_Sub_2_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_0__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_2_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_U3 ( .A(r[0]), 
        .B(r[1]), .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_3_), .B2(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[1]), .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_1__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[2]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_2_rs1[1]), .C2(Midori_rounds_sub_Sub_2_rs1[2]), 
        .A(Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_2_rs1[1]), .A2(Midori_rounds_sub_Sub_2_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_rs2[1]), .B(Midori_rounds_sub_Sub_2_rs2[0]), 
        .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_U1 ( .A(r[2]), .B(
        r[1]), .Z(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_3__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_rs2[0]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_3__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[3]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_3__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_3__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_3__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_3__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_2_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_U3 ( .A(r[2]), 
        .B(r[3]), .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[3]), .B2(
        Midori_rounds_sub_Sub_2_rs1[4]), .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_2_rs1[5]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_4__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[5]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_rs2[1]), .B(Midori_rounds_sub_Sub_2_rs2[0]), 
        .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_U1 ( .A(r[4]), .B(
        r[3]), .Z(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_6__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_rs2[0]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_6__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[6]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_6__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_rs1[4]), .C2(Midori_rounds_sub_Sub_2_rs1[5]), 
        .A(Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_6__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_6__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_rs1[4]), .A2(Midori_rounds_sub_Sub_2_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_6__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[7]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_2_rs1[4]), .C2(Midori_rounds_sub_Sub_2_rs1[5]), 
        .A(Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_rs1[4]), .A2(Midori_rounds_sub_Sub_2_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_2_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_U1 ( .A(r[4]), 
        .B(r[5]), .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_7__CF_Inst_n9) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_n21), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_n20), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[8]) );
  OAI21_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_U5 ( .B1(
        Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_3_), .B2(
        Midori_rounds_sub_Sub_2_rs1[1]), .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_n19), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_n20) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_2_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_n19) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_n18), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_n17), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_n21) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_rs2[1]), .B(r[5]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_n17) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_rs2[0]), .B(r[0]), .Z(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_8__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_9__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_rs2[2]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_9__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[9]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_9__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_rs1[1]), .C2(Midori_rounds_sub_Sub_2_rs1[2]), 
        .A(Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_9__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_9__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_rs1[1]), .A2(Midori_rounds_sub_Sub_2_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_9__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_U3 ( .A(r[6]), 
        .B(r[7]), .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[2]), .B1(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_10__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[11]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_2_rs1[1]), .C2(Midori_rounds_sub_Sub_2_rs1[2]), 
        .A(Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_2_rs1[1]), .A2(Midori_rounds_sub_Sub_2_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_rs2[3]), .B(Midori_rounds_sub_Sub_2_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_U1 ( .A(r[8]), 
        .B(r[7]), .Z(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_rs2[2]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[12]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_12__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_12__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_12__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_U3 ( .A(r[8]), 
        .B(r[9]), .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_2_rs1[5]), .B1(Midori_rounds_sub_Sub_2_rs1[4]), 
        .B2(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_13__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[14]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_rs2[3]), .B(Midori_rounds_sub_Sub_2_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_U1 ( .A(r[10]), 
        .B(r[9]), .Z(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_15__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_rs2[2]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_15__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[15]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_15__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_rs1[4]), .C2(Midori_rounds_sub_Sub_2_rs1[5]), 
        .A(Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_15__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_15__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_rs1[4]), .A2(Midori_rounds_sub_Sub_2_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_15__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[16]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_2_rs1[4]), .C2(Midori_rounds_sub_Sub_2_rs1[5]), 
        .A(Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_rs1[4]), .A2(Midori_rounds_sub_Sub_2_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_2_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_U1 ( .A(r[10]), 
        .B(r[11]), .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_16__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_U4 ( .A(r[6]), 
        .B(Midori_rounds_sub_Sub_2_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_n16) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_U3 ( .A(r[11]), 
        .B(Midori_rounds_sub_Sub_2_rs2[3]), .Z(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_n17) );
  AOI22_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_2_rs1[2]), .B1(Midori_rounds_sub_Sub_2_rs1[1]), 
        .B2(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_17__CF_Inst_n15) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_18__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_rs2[4]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_18__CF_Inst_n3), .Z(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_rs1[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_18__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_U2 ( .A(r[13]), 
        .B(r[12]), .Z(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_rs2[5]), .B(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_19__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_2_rs1[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_U4 ( .A(r[13]), 
        .B(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_U2 ( .A(r[14]), 
        .B(Midori_rounds_sub_Sub_2_rs1[0]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_rs2[4]), .B(Midori_rounds_sub_Sub_2_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_20__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_21__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_21__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_2_rs2[4]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[21]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_21__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_rs1[4]), .A2(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_U2 ( .A(r[15]), 
        .B(r[14]), .Z(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_rs2[5]), .B(Midori_rounds_sub_Sub_2_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_22__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[23]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_U4 ( .A(r[15]), 
        .B(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_U2 ( .A(r[16]), 
        .B(Midori_rounds_sub_Sub_2_S1_InAff_out3_reg[0]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_rs2[4]), .B(Midori_rounds_sub_Sub_2_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_23__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_24__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_24__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_2_rs2[4]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[24]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_rs1[4]), .A2(
        Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_24__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[25]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_rs1[4]), .A2(
        Midori_rounds_sub_Sub_2_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_U2 ( .A(r[17]), 
        .B(r[16]), .Z(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_rs2[5]), .B(Midori_rounds_sub_Sub_2_rs1[3]), 
        .ZN(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_2_rs1[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_U4 ( .A(r[17]), 
        .B(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_U2 ( .A(r[12]), 
        .B(Midori_rounds_sub_Sub_2_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_rs2[4]), .B(Midori_rounds_sub_Sub_2_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_2_S1_F_inst_Inst_26__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_1__Compression2_n2), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_1__Compression2_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_2_S1_F_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_2_S1_F_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[37]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result1[37]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[37]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_0__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_0__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[0]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_0__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_U2 ( .A(r[31]), 
        .B(r[30]), .Z(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_2_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_1__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_U2 ( .A(1'b0), .B(
        r[32]), .Z(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_U1 ( .A(1'b0), 
        .B(r[31]), .ZN(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_3__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_3__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_U2 ( .A(r[33]), 
        .B(r[32]), .Z(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_2_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_4__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[5]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_U2 ( .A(1'b0), .B(
        r[34]), .Z(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_U1 ( .A(1'b0), 
        .B(r[33]), .ZN(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_6__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_6__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[6]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_6__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_7__CF_Inst_U4 ( .A(1'b0), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_7__CF_Inst_n9), .Z(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_7__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_7__CF_Inst_n8), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_7__CF_Inst_n7), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_7__CF_Inst_n9) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_7__CF_Inst_n7) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_7__CF_Inst_U1 ( .A(r[34]), 
        .B(r[35]), .Z(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_7__CF_Inst_n8) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_U4 ( .A(r[35]), 
        .B(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_U2 ( .A(r[30]), 
        .B(Midori_rounds_sub_Sub_2_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_U1 ( .A(1'b0), .B(
        1'b0), .Z(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_8__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_9__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_9__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[9]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[1]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_U1 ( .A(r[18]), 
        .B(r[19]), .Z(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_10__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[11]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_U4 ( .A(r[19]), 
        .B(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_U2 ( .A(r[20]), 
        .B(Midori_rounds_sub_Sub_2_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_12__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[1]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_U1 ( .A(r[20]), 
        .B(r[21]), .Z(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_13__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[14]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_U4 ( .A(r[21]), 
        .B(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_U2 ( .A(r[22]), 
        .B(Midori_rounds_sub_Sub_2_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_15__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_15__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[15]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_U2 ( .A(r[23]), 
        .B(r[22]), .Z(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_2_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_n13), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_n12), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_n12) );
  INV_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[1]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_U2 ( .A(r[23]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_n13)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_U1 ( .A(r[18]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_17__CF_Inst_n15)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_18__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_18__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[18]) );
  AOI21_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_18__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_18__CF_Inst_n6) );
  OAI21_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_18__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_U3 ( .A(r[24]), 
        .B(r[25]), .ZN(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[2]), .B1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[1]), .B2(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_19__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[20]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[1]), .C2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_U1 ( .A(r[26]), 
        .B(r[25]), .Z(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_20__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_21__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_21__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[21]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_21__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_21__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_U3 ( .A(r[26]), 
        .B(r[27]), .ZN(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[2]), .B1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[1]), .B2(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_22__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[23]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_U1 ( .A(r[28]), 
        .B(r[27]), .Z(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_23__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_24__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_24__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[24]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_24__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[25]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[3]), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_n9), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_U1 ( .A(r[28]), 
        .B(r[29]), .ZN(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_25__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Out[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_U4 ( .A(r[24]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_n16)
         );
  XOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_U3 ( .A(r[29]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_n17)
         );
  AOI22_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[2]), .B1(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[36]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[36]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[36]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[38]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[38]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[38]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[39]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[39]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[39]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_2_S1_G_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_2_S1_G_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_InAff_out3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_S2_InAff_out3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_InAff_out3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_S2_InAff_out3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_InAff_out3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_S2_InAff_out3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_InAff_out3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_2_S2_InAff_out3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_S2_InAff_out2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_rs2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_S2_InAff_out2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_rs2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_S2_InAff_out2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_rs2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_2_S2_InAff_out2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_3_), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_S2_InAff_out1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_rs2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_S2_InAff_out1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_rs2[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_S2_InAff_out1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_rs2[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_2_S2_InAff_out1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_3_), .QN() );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_InputAffine_U3 ( .A(
        Midori_rounds_sub_Sub_2_S2_InAff_out3[1]), .B(Midori_rounds_n939), .Z(
        Midori_rounds_sub_Sub_2_S2_InAff_out3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_InputAffine_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_InAff_out2[1]), .B(Midori_rounds_n875), .Z(
        Midori_rounds_sub_Sub_2_S2_InAff_out2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_InputAffine_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_InAff_out1[1]), .B(Midori_rounds_n821), .Z(
        Midori_rounds_sub_Sub_2_S2_InAff_out1[3]) );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_rs2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_rs2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_0__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_rs1[0]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_0__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[0]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_0__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_rs2[1]), .C2(Midori_rounds_sub_Sub_2_rs2[2]), 
        .A(Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_0__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_0__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_rs2[1]), .A2(Midori_rounds_sub_Sub_2_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_0__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_2_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_U3 ( .A(r[36]), 
        .B(r[37]), .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_3_), .B2(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[1]), .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_1__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[2]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_2_rs2[1]), .C2(Midori_rounds_sub_Sub_2_rs2[2]), 
        .A(Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_2_rs2[1]), .A2(Midori_rounds_sub_Sub_2_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_rs1[1]), .B(Midori_rounds_sub_Sub_2_rs1[0]), 
        .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_U1 ( .A(r[38]), 
        .B(r[37]), .Z(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_3__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_rs1[0]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_3__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[3]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_3__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_3__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_3__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_3__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_2_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_U3 ( .A(r[38]), 
        .B(r[39]), .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[3]), .B2(
        Midori_rounds_sub_Sub_2_rs2[4]), .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_2_rs2[5]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_4__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[5]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_rs1[1]), .B(Midori_rounds_sub_Sub_2_rs1[0]), 
        .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_U1 ( .A(r[40]), 
        .B(r[39]), .Z(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_6__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_rs1[0]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_6__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[6]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_6__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_rs2[4]), .C2(Midori_rounds_sub_Sub_2_rs2[5]), 
        .A(Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_6__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_6__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_rs2[4]), .A2(Midori_rounds_sub_Sub_2_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_6__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[7]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_2_rs2[4]), .C2(Midori_rounds_sub_Sub_2_rs2[5]), 
        .A(Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_rs2[4]), .A2(Midori_rounds_sub_Sub_2_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_2_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_U1 ( .A(r[40]), 
        .B(r[41]), .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_7__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_n21), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_n20), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[8]) );
  OAI21_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_U5 ( .B1(
        Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_3_), .B2(
        Midori_rounds_sub_Sub_2_rs2[1]), .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_n19), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_n20) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_2_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_n19) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_n18), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_n17), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_n21) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_rs1[1]), .B(r[41]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_n17) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_rs1[0]), .B(r[36]), .Z(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_8__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_9__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_rs1[2]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_9__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[9]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_9__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_rs2[1]), .C2(Midori_rounds_sub_Sub_2_rs2[2]), 
        .A(Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_9__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_9__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_rs2[1]), .A2(Midori_rounds_sub_Sub_2_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_9__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_U3 ( .A(r[42]), 
        .B(r[43]), .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[2]), .B1(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[1]), .B2(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_10__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[11]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_2_rs2[1]), .C2(Midori_rounds_sub_Sub_2_rs2[2]), 
        .A(Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_2_rs2[1]), .A2(Midori_rounds_sub_Sub_2_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_rs1[3]), .B(Midori_rounds_sub_Sub_2_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_U1 ( .A(r[44]), 
        .B(r[43]), .Z(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_rs1[2]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[12]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_12__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_12__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_12__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_U3 ( .A(r[44]), 
        .B(r[45]), .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_2_rs2[5]), .B1(Midori_rounds_sub_Sub_2_rs2[4]), 
        .B2(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_13__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[14]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_rs1[3]), .B(Midori_rounds_sub_Sub_2_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_U1 ( .A(r[46]), 
        .B(r[45]), .Z(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_15__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_rs1[2]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_15__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[15]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_15__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_rs2[4]), .C2(Midori_rounds_sub_Sub_2_rs2[5]), 
        .A(Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_15__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_15__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_rs2[4]), .A2(Midori_rounds_sub_Sub_2_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_15__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[16]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_2_rs2[4]), .C2(Midori_rounds_sub_Sub_2_rs2[5]), 
        .A(Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_rs2[4]), .A2(Midori_rounds_sub_Sub_2_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_2_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_U1 ( .A(r[46]), 
        .B(r[47]), .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_16__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_U4 ( .A(r[42]), 
        .B(Midori_rounds_sub_Sub_2_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_n16) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_U3 ( .A(r[47]), 
        .B(Midori_rounds_sub_Sub_2_rs1[3]), .Z(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_n17) );
  AOI22_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_2_rs2[2]), .B1(Midori_rounds_sub_Sub_2_rs2[1]), 
        .B2(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_17__CF_Inst_n15) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_18__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_rs1[4]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_18__CF_Inst_n3), .Z(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_rs2[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_18__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_U2 ( .A(r[49]), 
        .B(r[48]), .Z(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_rs1[5]), .B(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_19__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_2_rs2[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_U4 ( .A(r[49]), 
        .B(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_U2 ( .A(r[50]), 
        .B(Midori_rounds_sub_Sub_2_rs2[0]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_rs1[4]), .B(Midori_rounds_sub_Sub_2_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_20__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_21__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_21__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_2_rs1[4]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[21]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_21__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_rs2[4]), .A2(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_U2 ( .A(r[51]), 
        .B(r[50]), .Z(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_rs1[5]), .B(Midori_rounds_sub_Sub_2_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_22__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[23]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_U4 ( .A(r[51]), 
        .B(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_U2 ( .A(r[52]), 
        .B(Midori_rounds_sub_Sub_2_S2_InAff_out3_reg[0]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_rs1[4]), .B(Midori_rounds_sub_Sub_2_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_23__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_24__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_24__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_2_rs1[4]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[24]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_rs2[4]), .A2(
        Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_24__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[25]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_rs2[4]), .A2(
        Midori_rounds_sub_Sub_2_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_U2 ( .A(r[53]), 
        .B(r[52]), .Z(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_rs1[5]), .B(Midori_rounds_sub_Sub_2_rs2[3]), 
        .ZN(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_2_rs2[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_U4 ( .A(r[53]), 
        .B(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_U2 ( .A(r[48]), 
        .B(Midori_rounds_sub_Sub_2_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_rs1[4]), .B(Midori_rounds_sub_Sub_2_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_2_S2_F_inst_Inst_26__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_1__Compression2_n2), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_1__Compression2_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_2_S2_F_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_2_S2_F_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[57]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result1[57]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[57]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_0__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_0__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[0]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_0__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_U2 ( .A(r[67]), 
        .B(r[66]), .Z(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_2_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_1__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_U2 ( .A(1'b0), .B(
        r[68]), .Z(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_U1 ( .A(1'b0), 
        .B(r[67]), .ZN(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_3__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_3__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_U2 ( .A(r[69]), 
        .B(r[68]), .Z(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_2_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_4__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[5]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_U2 ( .A(1'b0), .B(
        r[70]), .Z(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_U1 ( .A(1'b0), 
        .B(r[69]), .ZN(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_6__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_6__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[6]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_6__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_7__CF_Inst_U4 ( .A(1'b0), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_7__CF_Inst_n9), .Z(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_7__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_7__CF_Inst_n8), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_7__CF_Inst_n7), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_7__CF_Inst_n9) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_7__CF_Inst_n7) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_7__CF_Inst_U1 ( .A(r[70]), 
        .B(r[71]), .Z(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_7__CF_Inst_n8) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_U4 ( .A(r[71]), 
        .B(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_U2 ( .A(r[66]), 
        .B(Midori_rounds_sub_Sub_2_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_U1 ( .A(1'b0), .B(
        1'b0), .Z(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_8__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_9__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_9__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[9]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[1]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_U1 ( .A(r[54]), 
        .B(r[55]), .Z(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_10__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[11]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_U4 ( .A(r[55]), 
        .B(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_U2 ( .A(r[56]), 
        .B(Midori_rounds_sub_Sub_2_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_12__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[1]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_U1 ( .A(r[56]), 
        .B(r[57]), .Z(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_13__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[14]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_U4 ( .A(r[57]), 
        .B(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_U2 ( .A(r[58]), 
        .B(Midori_rounds_sub_Sub_2_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_15__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_15__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[15]) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_U2 ( .A(r[59]), 
        .B(r[58]), .Z(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_2_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_n13), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_n12), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_n12) );
  INV_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[1]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_U2 ( .A(r[59]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_n13)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_U1 ( .A(r[54]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_17__CF_Inst_n15)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_18__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_18__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[18]) );
  AOI21_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_18__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_18__CF_Inst_n6) );
  OAI21_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_18__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_U3 ( .A(r[60]), 
        .B(r[61]), .ZN(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[2]), .B1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[1]), .B2(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_19__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[20]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[1]), .C2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_U1 ( .A(r[62]), 
        .B(r[61]), .Z(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_20__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_21__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_21__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[21]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_21__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_21__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_U3 ( .A(r[62]), 
        .B(r[63]), .ZN(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[2]), .B1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[1]), .B2(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_22__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[23]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_U1 ( .A(r[64]), 
        .B(r[63]), .Z(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_23__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_24__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_24__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[24]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_24__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[25]) );
  OAI211_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[3]), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_n9), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_U1 ( .A(r[64]), 
        .B(r[65]), .ZN(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_25__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Out[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_U4 ( .A(r[60]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_n16)
         );
  XOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_U3 ( .A(r[65]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_n17)
         );
  AOI22_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[2]), .B1(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[56]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[56]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[56]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[58]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[58]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[58]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[59]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[59]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[59]) );
  XNOR2_X1 Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_2_S2_G_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_2_S2_G_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_InAff_out3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_S1_InAff_out3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_InAff_out3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_S1_InAff_out3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_InAff_out3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_S1_InAff_out3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_InAff_out3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_3_S1_InAff_out3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_S1_InAff_out2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_rs1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_S1_InAff_out2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_rs1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_S1_InAff_out2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_rs1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_3_S1_InAff_out2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_3_), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_S1_InAff_out1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_rs1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_S1_InAff_out1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_rs1[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_S1_InAff_out1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_rs1[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_3_S1_InAff_out1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_3_), .QN() );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_InputAffine_U3 ( .A(
        Midori_rounds_sub_Sub_3_S1_InAff_out3[1]), .B(Midori_rounds_n943), .Z(
        Midori_rounds_sub_Sub_3_S1_InAff_out3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_InputAffine_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_InAff_out2[1]), .B(Midori_rounds_n879), .Z(
        Midori_rounds_sub_Sub_3_S1_InAff_out2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_InputAffine_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_InAff_out1[1]), .B(Midori_rounds_n824), .Z(
        Midori_rounds_sub_Sub_3_S1_InAff_out1[3]) );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_rs1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_rs1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_0__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_rs2[0]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_0__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[0]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_0__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_rs1[1]), .C2(Midori_rounds_sub_Sub_3_rs1[2]), 
        .A(Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_0__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_0__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_rs1[1]), .A2(Midori_rounds_sub_Sub_3_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_0__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_3_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_U3 ( .A(r[0]), 
        .B(r[1]), .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_3_), .B2(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[1]), .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_1__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[2]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_3_rs1[1]), .C2(Midori_rounds_sub_Sub_3_rs1[2]), 
        .A(Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_3_rs1[1]), .A2(Midori_rounds_sub_Sub_3_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_rs2[1]), .B(Midori_rounds_sub_Sub_3_rs2[0]), 
        .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_U1 ( .A(r[2]), .B(
        r[1]), .Z(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_3__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_rs2[0]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_3__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[3]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_3__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_3__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_3__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_3__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_3_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_U3 ( .A(r[2]), 
        .B(r[3]), .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[3]), .B2(
        Midori_rounds_sub_Sub_3_rs1[4]), .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_3_rs1[5]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_4__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[5]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_rs2[1]), .B(Midori_rounds_sub_Sub_3_rs2[0]), 
        .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_U1 ( .A(r[4]), .B(
        r[3]), .Z(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_6__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_rs2[0]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_6__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[6]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_6__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_rs1[4]), .C2(Midori_rounds_sub_Sub_3_rs1[5]), 
        .A(Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_6__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_6__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_rs1[4]), .A2(Midori_rounds_sub_Sub_3_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_6__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[7]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_3_rs1[4]), .C2(Midori_rounds_sub_Sub_3_rs1[5]), 
        .A(Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_rs1[4]), .A2(Midori_rounds_sub_Sub_3_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_3_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_U1 ( .A(r[4]), 
        .B(r[5]), .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_7__CF_Inst_n9) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_n21), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_n20), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[8]) );
  OAI21_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_U5 ( .B1(
        Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_3_), .B2(
        Midori_rounds_sub_Sub_3_rs1[1]), .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_n19), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_n20) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_3_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_n19) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_n18), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_n17), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_n21) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_rs2[1]), .B(r[5]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_n17) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_rs2[0]), .B(r[0]), .Z(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_8__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_9__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_rs2[2]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_9__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[9]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_9__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_rs1[1]), .C2(Midori_rounds_sub_Sub_3_rs1[2]), 
        .A(Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_9__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_9__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_rs1[1]), .A2(Midori_rounds_sub_Sub_3_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_9__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_U3 ( .A(r[6]), 
        .B(r[7]), .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[2]), .B1(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_10__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[11]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_3_rs1[1]), .C2(Midori_rounds_sub_Sub_3_rs1[2]), 
        .A(Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_3_rs1[1]), .A2(Midori_rounds_sub_Sub_3_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_rs2[3]), .B(Midori_rounds_sub_Sub_3_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_U1 ( .A(r[8]), 
        .B(r[7]), .Z(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_rs2[2]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[12]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_12__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_12__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_12__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_U3 ( .A(r[8]), 
        .B(r[9]), .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_3_rs1[5]), .B1(Midori_rounds_sub_Sub_3_rs1[4]), 
        .B2(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_13__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[14]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_rs2[3]), .B(Midori_rounds_sub_Sub_3_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_U1 ( .A(r[10]), 
        .B(r[9]), .Z(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_15__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_rs2[2]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_15__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[15]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_15__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_rs1[4]), .C2(Midori_rounds_sub_Sub_3_rs1[5]), 
        .A(Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_15__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_15__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_rs1[4]), .A2(Midori_rounds_sub_Sub_3_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_15__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[16]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_3_rs1[4]), .C2(Midori_rounds_sub_Sub_3_rs1[5]), 
        .A(Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_rs1[4]), .A2(Midori_rounds_sub_Sub_3_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_3_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_U1 ( .A(r[10]), 
        .B(r[11]), .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_16__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_U4 ( .A(r[6]), 
        .B(Midori_rounds_sub_Sub_3_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_n16) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_U3 ( .A(r[11]), 
        .B(Midori_rounds_sub_Sub_3_rs2[3]), .Z(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_n17) );
  AOI22_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_3_rs1[2]), .B1(Midori_rounds_sub_Sub_3_rs1[1]), 
        .B2(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_17__CF_Inst_n15) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_18__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_rs2[4]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_18__CF_Inst_n3), .Z(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_rs1[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_18__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_U2 ( .A(r[13]), 
        .B(r[12]), .Z(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_rs2[5]), .B(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_19__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_3_rs1[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_U4 ( .A(r[13]), 
        .B(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_U2 ( .A(r[14]), 
        .B(Midori_rounds_sub_Sub_3_rs1[0]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_rs2[4]), .B(Midori_rounds_sub_Sub_3_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_20__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_21__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_21__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_3_rs2[4]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[21]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_21__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_rs1[4]), .A2(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_U2 ( .A(r[15]), 
        .B(r[14]), .Z(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_rs2[5]), .B(Midori_rounds_sub_Sub_3_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_22__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[23]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_U4 ( .A(r[15]), 
        .B(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_U2 ( .A(r[16]), 
        .B(Midori_rounds_sub_Sub_3_S1_InAff_out3_reg[0]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_rs2[4]), .B(Midori_rounds_sub_Sub_3_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_23__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_24__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_24__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_3_rs2[4]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[24]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_rs1[4]), .A2(
        Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_24__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[25]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_rs1[4]), .A2(
        Midori_rounds_sub_Sub_3_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_U2 ( .A(r[17]), 
        .B(r[16]), .Z(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_rs2[5]), .B(Midori_rounds_sub_Sub_3_rs1[3]), 
        .ZN(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_3_rs1[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_U4 ( .A(r[17]), 
        .B(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_U2 ( .A(r[12]), 
        .B(Midori_rounds_sub_Sub_3_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_rs2[4]), .B(Midori_rounds_sub_Sub_3_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_3_S1_F_inst_Inst_26__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_1__Compression2_n2), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_1__Compression2_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_3_S1_F_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_3_S1_F_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result1[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[29]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_0__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_0__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[0]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_0__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_U2 ( .A(r[31]), 
        .B(r[30]), .Z(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_3_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_1__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_U2 ( .A(1'b0), .B(
        r[32]), .Z(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_U1 ( .A(1'b0), 
        .B(r[31]), .ZN(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_3__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_3__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_U2 ( .A(r[33]), 
        .B(r[32]), .Z(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_3_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_4__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[5]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_U2 ( .A(1'b0), .B(
        r[34]), .Z(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_U1 ( .A(1'b0), 
        .B(r[33]), .ZN(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_6__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_6__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[6]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_6__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_7__CF_Inst_U4 ( .A(1'b0), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_7__CF_Inst_n9), .Z(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_7__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_7__CF_Inst_n8), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_7__CF_Inst_n7), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_7__CF_Inst_n9) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_7__CF_Inst_n7) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_7__CF_Inst_U1 ( .A(r[34]), 
        .B(r[35]), .Z(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_7__CF_Inst_n8) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_U4 ( .A(r[35]), 
        .B(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_U2 ( .A(r[30]), 
        .B(Midori_rounds_sub_Sub_3_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_U1 ( .A(1'b0), .B(
        1'b0), .Z(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_8__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_9__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_9__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[9]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[1]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_U1 ( .A(r[18]), 
        .B(r[19]), .Z(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_10__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[11]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_U4 ( .A(r[19]), 
        .B(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_U2 ( .A(r[20]), 
        .B(Midori_rounds_sub_Sub_3_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_12__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[1]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_U1 ( .A(r[20]), 
        .B(r[21]), .Z(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_13__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[14]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_U4 ( .A(r[21]), 
        .B(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_U2 ( .A(r[22]), 
        .B(Midori_rounds_sub_Sub_3_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_15__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_15__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[15]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_U2 ( .A(r[23]), 
        .B(r[22]), .Z(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_3_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_n13), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_n12), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_n12) );
  INV_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[1]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_U2 ( .A(r[23]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_n13)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_U1 ( .A(r[18]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_17__CF_Inst_n15)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_18__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_18__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[18]) );
  AOI21_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_18__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_18__CF_Inst_n6) );
  OAI21_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_18__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_U3 ( .A(r[24]), 
        .B(r[25]), .ZN(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[2]), .B1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[1]), .B2(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_19__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[20]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[1]), .C2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_U1 ( .A(r[26]), 
        .B(r[25]), .Z(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_20__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_21__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_21__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[21]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_21__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_21__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_U3 ( .A(r[26]), 
        .B(r[27]), .ZN(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[2]), .B1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[1]), .B2(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_22__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[23]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_U1 ( .A(r[28]), 
        .B(r[27]), .Z(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_23__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_24__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_24__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[24]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_24__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[25]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[3]), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_n9), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_U1 ( .A(r[28]), 
        .B(r[29]), .ZN(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_25__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Out[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_U4 ( .A(r[24]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_n16)
         );
  XOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_U3 ( .A(r[29]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_n17)
         );
  AOI22_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[2]), .B1(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[28]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[28]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[28]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[30]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[30]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[30]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[31]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[31]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[31]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_3_S1_G_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_3_S1_G_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_InAff_out3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_S2_InAff_out3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_InAff_out3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_S2_InAff_out3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_InAff_out3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_S2_InAff_out3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_InAff_out3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_3_S2_InAff_out3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_S2_InAff_out2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_rs2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_S2_InAff_out2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_rs2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_S2_InAff_out2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_rs2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_3_S2_InAff_out2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_3_), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_S2_InAff_out1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_rs2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_S2_InAff_out1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_rs2[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_S2_InAff_out1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_rs2[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_3_S2_InAff_out1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_3_), .QN() );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_InputAffine_U3 ( .A(
        Midori_rounds_sub_Sub_3_S2_InAff_out3[1]), .B(Midori_rounds_n947), .Z(
        Midori_rounds_sub_Sub_3_S2_InAff_out3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_InputAffine_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_InAff_out2[1]), .B(Midori_rounds_n883), .Z(
        Midori_rounds_sub_Sub_3_S2_InAff_out2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_InputAffine_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_InAff_out1[1]), .B(Midori_rounds_n827), .Z(
        Midori_rounds_sub_Sub_3_S2_InAff_out1[3]) );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_rs2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_rs2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_0__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_rs1[0]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_0__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[0]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_0__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_rs2[1]), .C2(Midori_rounds_sub_Sub_3_rs2[2]), 
        .A(Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_0__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_0__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_rs2[1]), .A2(Midori_rounds_sub_Sub_3_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_0__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_3_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_U3 ( .A(r[36]), 
        .B(r[37]), .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_3_), .B2(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[1]), .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_1__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[2]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_3_rs2[1]), .C2(Midori_rounds_sub_Sub_3_rs2[2]), 
        .A(Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_3_rs2[1]), .A2(Midori_rounds_sub_Sub_3_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_rs1[1]), .B(Midori_rounds_sub_Sub_3_rs1[0]), 
        .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_U1 ( .A(r[38]), 
        .B(r[37]), .Z(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_3__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_rs1[0]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_3__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[3]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_3__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_3__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_3__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_3__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_3_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_U3 ( .A(r[38]), 
        .B(r[39]), .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[3]), .B2(
        Midori_rounds_sub_Sub_3_rs2[4]), .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_3_rs2[5]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_4__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[5]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_rs1[1]), .B(Midori_rounds_sub_Sub_3_rs1[0]), 
        .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_U1 ( .A(r[40]), 
        .B(r[39]), .Z(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_6__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_rs1[0]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_6__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[6]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_6__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_rs2[4]), .C2(Midori_rounds_sub_Sub_3_rs2[5]), 
        .A(Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_6__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_6__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_rs2[4]), .A2(Midori_rounds_sub_Sub_3_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_6__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[7]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_3_rs2[4]), .C2(Midori_rounds_sub_Sub_3_rs2[5]), 
        .A(Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_rs2[4]), .A2(Midori_rounds_sub_Sub_3_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_3_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_U1 ( .A(r[40]), 
        .B(r[41]), .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_7__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_n21), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_n20), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[8]) );
  OAI21_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_U5 ( .B1(
        Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_3_), .B2(
        Midori_rounds_sub_Sub_3_rs2[1]), .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_n19), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_n20) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_3_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_n19) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_n18), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_n17), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_n21) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_rs1[1]), .B(r[41]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_n17) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_rs1[0]), .B(r[36]), .Z(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_8__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_9__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_rs1[2]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_9__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[9]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_9__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_rs2[1]), .C2(Midori_rounds_sub_Sub_3_rs2[2]), 
        .A(Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_9__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_9__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_rs2[1]), .A2(Midori_rounds_sub_Sub_3_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_9__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_U3 ( .A(r[42]), 
        .B(r[43]), .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[2]), .B1(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[1]), .B2(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_10__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[11]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_3_rs2[1]), .C2(Midori_rounds_sub_Sub_3_rs2[2]), 
        .A(Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_3_rs2[1]), .A2(Midori_rounds_sub_Sub_3_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_rs1[3]), .B(Midori_rounds_sub_Sub_3_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_U1 ( .A(r[44]), 
        .B(r[43]), .Z(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_rs1[2]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[12]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_12__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_12__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_12__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_U3 ( .A(r[44]), 
        .B(r[45]), .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_3_rs2[5]), .B1(Midori_rounds_sub_Sub_3_rs2[4]), 
        .B2(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_13__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[14]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_rs1[3]), .B(Midori_rounds_sub_Sub_3_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_U1 ( .A(r[46]), 
        .B(r[45]), .Z(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_15__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_rs1[2]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_15__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[15]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_15__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_rs2[4]), .C2(Midori_rounds_sub_Sub_3_rs2[5]), 
        .A(Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_15__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_15__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_rs2[4]), .A2(Midori_rounds_sub_Sub_3_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_15__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[16]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_3_rs2[4]), .C2(Midori_rounds_sub_Sub_3_rs2[5]), 
        .A(Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_rs2[4]), .A2(Midori_rounds_sub_Sub_3_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_3_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_U1 ( .A(r[46]), 
        .B(r[47]), .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_16__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_U4 ( .A(r[42]), 
        .B(Midori_rounds_sub_Sub_3_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_n16) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_U3 ( .A(r[47]), 
        .B(Midori_rounds_sub_Sub_3_rs1[3]), .Z(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_n17) );
  AOI22_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_3_rs2[2]), .B1(Midori_rounds_sub_Sub_3_rs2[1]), 
        .B2(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_17__CF_Inst_n15) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_18__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_rs1[4]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_18__CF_Inst_n3), .Z(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_rs2[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_18__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_U2 ( .A(r[49]), 
        .B(r[48]), .Z(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_rs1[5]), .B(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_19__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_3_rs2[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_U4 ( .A(r[49]), 
        .B(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_U2 ( .A(r[50]), 
        .B(Midori_rounds_sub_Sub_3_rs2[0]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_rs1[4]), .B(Midori_rounds_sub_Sub_3_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_20__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_21__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_21__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_3_rs1[4]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[21]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_21__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_rs2[4]), .A2(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_U2 ( .A(r[51]), 
        .B(r[50]), .Z(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_rs1[5]), .B(Midori_rounds_sub_Sub_3_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_22__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[23]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_U4 ( .A(r[51]), 
        .B(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_U2 ( .A(r[52]), 
        .B(Midori_rounds_sub_Sub_3_S2_InAff_out3_reg[0]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_rs1[4]), .B(Midori_rounds_sub_Sub_3_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_23__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_24__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_24__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_3_rs1[4]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[24]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_rs2[4]), .A2(
        Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_24__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[25]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_rs2[4]), .A2(
        Midori_rounds_sub_Sub_3_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_U2 ( .A(r[53]), 
        .B(r[52]), .Z(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_rs1[5]), .B(Midori_rounds_sub_Sub_3_rs2[3]), 
        .ZN(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_3_rs2[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_U4 ( .A(r[53]), 
        .B(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_U2 ( .A(r[48]), 
        .B(Midori_rounds_sub_Sub_3_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_rs1[4]), .B(Midori_rounds_sub_Sub_3_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_3_S2_F_inst_Inst_26__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_1__Compression2_n2), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_1__Compression2_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_3_S2_F_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_3_S2_F_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_0__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_0__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[0]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_0__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_U2 ( .A(r[67]), 
        .B(r[66]), .Z(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_3_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_1__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_U2 ( .A(1'b0), .B(
        r[68]), .Z(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_U1 ( .A(1'b0), 
        .B(r[67]), .ZN(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_3__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_3__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_U2 ( .A(r[69]), 
        .B(r[68]), .Z(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_3_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_4__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[5]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_U2 ( .A(1'b0), .B(
        r[70]), .Z(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_U1 ( .A(1'b0), 
        .B(r[69]), .ZN(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_6__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_6__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[6]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_6__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_7__CF_Inst_U4 ( .A(1'b0), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_7__CF_Inst_n9), .Z(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_7__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_7__CF_Inst_n8), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_7__CF_Inst_n7), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_7__CF_Inst_n9) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_7__CF_Inst_n7) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_7__CF_Inst_U1 ( .A(r[70]), 
        .B(r[71]), .Z(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_7__CF_Inst_n8) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_U4 ( .A(r[71]), 
        .B(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_U2 ( .A(r[66]), 
        .B(Midori_rounds_sub_Sub_3_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_U1 ( .A(1'b0), .B(
        1'b0), .Z(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_8__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_9__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_9__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[9]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[1]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_U1 ( .A(r[54]), 
        .B(r[55]), .Z(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_10__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[11]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_U4 ( .A(r[55]), 
        .B(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_U2 ( .A(r[56]), 
        .B(Midori_rounds_sub_Sub_3_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_12__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[1]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_U1 ( .A(r[56]), 
        .B(r[57]), .Z(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_13__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[14]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_U4 ( .A(r[57]), 
        .B(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_U2 ( .A(r[58]), 
        .B(Midori_rounds_sub_Sub_3_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_15__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_15__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[15]) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_U2 ( .A(r[59]), 
        .B(r[58]), .Z(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_3_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_n13), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_n12), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_n12) );
  INV_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[1]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_U2 ( .A(r[59]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_n13)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_U1 ( .A(r[54]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_17__CF_Inst_n15)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_18__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_18__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[18]) );
  AOI21_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_18__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_18__CF_Inst_n6) );
  OAI21_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_18__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_U3 ( .A(r[60]), 
        .B(r[61]), .ZN(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[2]), .B1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[1]), .B2(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_19__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[20]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[1]), .C2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_U1 ( .A(r[62]), 
        .B(r[61]), .Z(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_20__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_21__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_21__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[21]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_21__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_21__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_U3 ( .A(r[62]), 
        .B(r[63]), .ZN(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[2]), .B1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[1]), .B2(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_22__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[23]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_U1 ( .A(r[64]), 
        .B(r[63]), .Z(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_23__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_24__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_24__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[24]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_24__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[25]) );
  OAI211_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[3]), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_n9), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_U1 ( .A(r[64]), 
        .B(r[65]), .ZN(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_25__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Out[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_U4 ( .A(r[60]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_n16)
         );
  XOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_U3 ( .A(r[65]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_n17)
         );
  AOI22_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[2]), .B1(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_3_S2_G_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_3_S2_G_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_InAff_out3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_S1_InAff_out3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_InAff_out3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_S1_InAff_out3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_InAff_out3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_S1_InAff_out3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_InAff_out3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_4_S1_InAff_out3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_S1_InAff_out2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_rs1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_S1_InAff_out2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_rs1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_S1_InAff_out2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_rs1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_4_S1_InAff_out2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_3_), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_S1_InAff_out1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_rs1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_S1_InAff_out1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_rs1[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_S1_InAff_out1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_rs1[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_4_S1_InAff_out1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_3_), .QN() );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_InputAffine_U3 ( .A(
        Midori_rounds_sub_Sub_4_S1_InAff_out3[1]), .B(Midori_rounds_n951), .Z(
        Midori_rounds_sub_Sub_4_S1_InAff_out3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_InputAffine_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_InAff_out2[1]), .B(Midori_rounds_n887), .Z(
        Midori_rounds_sub_Sub_4_S1_InAff_out2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_InputAffine_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_InAff_out1[1]), .B(Midori_rounds_n830), .Z(
        Midori_rounds_sub_Sub_4_S1_InAff_out1[3]) );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_rs1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_rs1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_0__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_rs2[0]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_0__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[0]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_0__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_rs1[1]), .C2(Midori_rounds_sub_Sub_4_rs1[2]), 
        .A(Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_0__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_0__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_rs1[1]), .A2(Midori_rounds_sub_Sub_4_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_0__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_4_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_U3 ( .A(r[0]), 
        .B(r[1]), .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_3_), .B2(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[1]), .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_1__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[2]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_4_rs1[1]), .C2(Midori_rounds_sub_Sub_4_rs1[2]), 
        .A(Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_4_rs1[1]), .A2(Midori_rounds_sub_Sub_4_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_rs2[1]), .B(Midori_rounds_sub_Sub_4_rs2[0]), 
        .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_U1 ( .A(r[2]), .B(
        r[1]), .Z(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_3__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_rs2[0]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_3__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[3]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_3__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_3__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_3__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_3__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_4_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_U3 ( .A(r[2]), 
        .B(r[3]), .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[3]), .B2(
        Midori_rounds_sub_Sub_4_rs1[4]), .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_4_rs1[5]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_4__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[5]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_rs2[1]), .B(Midori_rounds_sub_Sub_4_rs2[0]), 
        .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_U1 ( .A(r[4]), .B(
        r[3]), .Z(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_6__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_rs2[0]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_6__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[6]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_6__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_rs1[4]), .C2(Midori_rounds_sub_Sub_4_rs1[5]), 
        .A(Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_6__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_6__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_rs1[4]), .A2(Midori_rounds_sub_Sub_4_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_6__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[7]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_4_rs1[4]), .C2(Midori_rounds_sub_Sub_4_rs1[5]), 
        .A(Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_rs1[4]), .A2(Midori_rounds_sub_Sub_4_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_4_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_U1 ( .A(r[4]), 
        .B(r[5]), .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_7__CF_Inst_n9) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_n21), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_n20), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[8]) );
  OAI21_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_U5 ( .B1(
        Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_3_), .B2(
        Midori_rounds_sub_Sub_4_rs1[1]), .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_n19), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_n20) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_4_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_n19) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_n18), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_n17), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_n21) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_rs2[1]), .B(r[5]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_n17) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_rs2[0]), .B(r[0]), .Z(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_8__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_9__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_rs2[2]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_9__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[9]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_9__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_rs1[1]), .C2(Midori_rounds_sub_Sub_4_rs1[2]), 
        .A(Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_9__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_9__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_rs1[1]), .A2(Midori_rounds_sub_Sub_4_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_9__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_U3 ( .A(r[6]), 
        .B(r[7]), .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[2]), .B1(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_10__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[11]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_4_rs1[1]), .C2(Midori_rounds_sub_Sub_4_rs1[2]), 
        .A(Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_4_rs1[1]), .A2(Midori_rounds_sub_Sub_4_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_rs2[3]), .B(Midori_rounds_sub_Sub_4_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_U1 ( .A(r[8]), 
        .B(r[7]), .Z(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_rs2[2]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[12]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_12__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_12__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_12__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_U3 ( .A(r[8]), 
        .B(r[9]), .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_4_rs1[5]), .B1(Midori_rounds_sub_Sub_4_rs1[4]), 
        .B2(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_13__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[14]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_rs2[3]), .B(Midori_rounds_sub_Sub_4_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_U1 ( .A(r[10]), 
        .B(r[9]), .Z(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_15__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_rs2[2]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_15__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[15]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_15__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_rs1[4]), .C2(Midori_rounds_sub_Sub_4_rs1[5]), 
        .A(Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_15__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_15__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_rs1[4]), .A2(Midori_rounds_sub_Sub_4_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_15__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[16]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_4_rs1[4]), .C2(Midori_rounds_sub_Sub_4_rs1[5]), 
        .A(Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_rs1[4]), .A2(Midori_rounds_sub_Sub_4_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_4_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_U1 ( .A(r[10]), 
        .B(r[11]), .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_16__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_U4 ( .A(r[6]), 
        .B(Midori_rounds_sub_Sub_4_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_n16) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_U3 ( .A(r[11]), 
        .B(Midori_rounds_sub_Sub_4_rs2[3]), .Z(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_n17) );
  AOI22_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_4_rs1[2]), .B1(Midori_rounds_sub_Sub_4_rs1[1]), 
        .B2(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_17__CF_Inst_n15) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_18__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_rs2[4]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_18__CF_Inst_n3), .Z(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_rs1[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_18__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_U2 ( .A(r[13]), 
        .B(r[12]), .Z(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_rs2[5]), .B(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_19__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_4_rs1[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_U4 ( .A(r[13]), 
        .B(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_U2 ( .A(r[14]), 
        .B(Midori_rounds_sub_Sub_4_rs1[0]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_rs2[4]), .B(Midori_rounds_sub_Sub_4_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_20__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_21__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_21__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_4_rs2[4]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[21]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_21__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_rs1[4]), .A2(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_U2 ( .A(r[15]), 
        .B(r[14]), .Z(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_rs2[5]), .B(Midori_rounds_sub_Sub_4_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_22__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[23]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_U4 ( .A(r[15]), 
        .B(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_U2 ( .A(r[16]), 
        .B(Midori_rounds_sub_Sub_4_S1_InAff_out3_reg[0]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_rs2[4]), .B(Midori_rounds_sub_Sub_4_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_23__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_24__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_24__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_4_rs2[4]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[24]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_rs1[4]), .A2(
        Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_24__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[25]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_rs1[4]), .A2(
        Midori_rounds_sub_Sub_4_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_U2 ( .A(r[17]), 
        .B(r[16]), .Z(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_rs2[5]), .B(Midori_rounds_sub_Sub_4_rs1[3]), 
        .ZN(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_4_rs1[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_U4 ( .A(r[17]), 
        .B(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_U2 ( .A(r[12]), 
        .B(Midori_rounds_sub_Sub_4_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_rs2[4]), .B(Midori_rounds_sub_Sub_4_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_4_S1_F_inst_Inst_26__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_1__Compression2_n2), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_1__Compression2_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_4_S1_F_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_4_S1_F_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result1[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_0__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_0__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[0]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_0__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_U2 ( .A(r[31]), 
        .B(r[30]), .Z(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_4_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_1__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_U2 ( .A(1'b0), .B(
        r[32]), .Z(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_U1 ( .A(1'b0), 
        .B(r[31]), .ZN(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_3__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_3__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_U2 ( .A(r[33]), 
        .B(r[32]), .Z(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_4_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_4__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[5]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_U2 ( .A(1'b0), .B(
        r[34]), .Z(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_U1 ( .A(1'b0), 
        .B(r[33]), .ZN(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_6__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_6__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[6]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_6__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_7__CF_Inst_U4 ( .A(1'b0), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_7__CF_Inst_n9), .Z(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_7__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_7__CF_Inst_n8), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_7__CF_Inst_n7), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_7__CF_Inst_n9) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_7__CF_Inst_n7) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_7__CF_Inst_U1 ( .A(r[34]), 
        .B(r[35]), .Z(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_7__CF_Inst_n8) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_U4 ( .A(r[35]), 
        .B(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_U2 ( .A(r[30]), 
        .B(Midori_rounds_sub_Sub_4_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_U1 ( .A(1'b0), .B(
        1'b0), .Z(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_8__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_9__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_9__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[9]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[1]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_U1 ( .A(r[18]), 
        .B(r[19]), .Z(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_10__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[11]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_U4 ( .A(r[19]), 
        .B(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_U2 ( .A(r[20]), 
        .B(Midori_rounds_sub_Sub_4_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_12__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[1]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_U1 ( .A(r[20]), 
        .B(r[21]), .Z(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_13__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[14]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_U4 ( .A(r[21]), 
        .B(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_U2 ( .A(r[22]), 
        .B(Midori_rounds_sub_Sub_4_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_15__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_15__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[15]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_U2 ( .A(r[23]), 
        .B(r[22]), .Z(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_4_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_n13), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_n12), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_n12) );
  INV_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[1]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_U2 ( .A(r[23]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_n13)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_U1 ( .A(r[18]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_17__CF_Inst_n15)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_18__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_18__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[18]) );
  AOI21_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_18__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_18__CF_Inst_n6) );
  OAI21_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_18__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_U3 ( .A(r[24]), 
        .B(r[25]), .ZN(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[2]), .B1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[1]), .B2(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_19__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[20]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[1]), .C2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_U1 ( .A(r[26]), 
        .B(r[25]), .Z(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_20__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_21__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_21__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[21]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_21__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_21__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_U3 ( .A(r[26]), 
        .B(r[27]), .ZN(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[2]), .B1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[1]), .B2(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_22__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[23]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_U1 ( .A(r[28]), 
        .B(r[27]), .Z(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_23__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_24__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_24__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[24]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_24__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[25]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[3]), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_n9), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_U1 ( .A(r[28]), 
        .B(r[29]), .ZN(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_25__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Out[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_U4 ( .A(r[24]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_n16)
         );
  XOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_U3 ( .A(r[29]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_n17)
         );
  AOI22_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[2]), .B1(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[12]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[12]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[12]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[14]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[14]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[14]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[15]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[15]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[15]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_4_S1_G_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_4_S1_G_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_InAff_out3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_S2_InAff_out3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_InAff_out3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_S2_InAff_out3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_InAff_out3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_S2_InAff_out3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_InAff_out3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_4_S2_InAff_out3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_S2_InAff_out2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_rs2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_S2_InAff_out2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_rs2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_S2_InAff_out2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_rs2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_4_S2_InAff_out2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_3_), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_S2_InAff_out1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_rs2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_S2_InAff_out1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_rs2[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_S2_InAff_out1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_rs2[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_4_S2_InAff_out1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_3_), .QN() );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_InputAffine_U3 ( .A(
        Midori_rounds_sub_Sub_4_S2_InAff_out3[1]), .B(Midori_rounds_n955), .Z(
        Midori_rounds_sub_Sub_4_S2_InAff_out3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_InputAffine_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_InAff_out2[1]), .B(Midori_rounds_n891), .Z(
        Midori_rounds_sub_Sub_4_S2_InAff_out2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_InputAffine_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_InAff_out1[1]), .B(Midori_rounds_n833), .Z(
        Midori_rounds_sub_Sub_4_S2_InAff_out1[3]) );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_rs2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_rs2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_0__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_rs1[0]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_0__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[0]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_0__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_rs2[1]), .C2(Midori_rounds_sub_Sub_4_rs2[2]), 
        .A(Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_0__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_0__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_rs2[1]), .A2(Midori_rounds_sub_Sub_4_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_0__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_4_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_U3 ( .A(r[36]), 
        .B(r[37]), .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_3_), .B2(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[1]), .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_1__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[2]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_4_rs2[1]), .C2(Midori_rounds_sub_Sub_4_rs2[2]), 
        .A(Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_4_rs2[1]), .A2(Midori_rounds_sub_Sub_4_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_rs1[1]), .B(Midori_rounds_sub_Sub_4_rs1[0]), 
        .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_U1 ( .A(r[38]), 
        .B(r[37]), .Z(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_3__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_rs1[0]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_3__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[3]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_3__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_3__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_3__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_3__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_4_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_U3 ( .A(r[38]), 
        .B(r[39]), .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[3]), .B2(
        Midori_rounds_sub_Sub_4_rs2[4]), .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_4_rs2[5]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_4__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[5]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_rs1[1]), .B(Midori_rounds_sub_Sub_4_rs1[0]), 
        .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_U1 ( .A(r[40]), 
        .B(r[39]), .Z(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_6__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_rs1[0]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_6__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[6]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_6__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_rs2[4]), .C2(Midori_rounds_sub_Sub_4_rs2[5]), 
        .A(Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_6__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_6__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_rs2[4]), .A2(Midori_rounds_sub_Sub_4_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_6__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[7]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_4_rs2[4]), .C2(Midori_rounds_sub_Sub_4_rs2[5]), 
        .A(Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_rs2[4]), .A2(Midori_rounds_sub_Sub_4_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_4_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_U1 ( .A(r[40]), 
        .B(r[41]), .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_7__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_n21), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_n20), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[8]) );
  OAI21_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_U5 ( .B1(
        Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_3_), .B2(
        Midori_rounds_sub_Sub_4_rs2[1]), .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_n19), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_n20) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_4_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_n19) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_n18), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_n17), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_n21) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_rs1[1]), .B(r[41]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_n17) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_rs1[0]), .B(r[36]), .Z(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_8__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_9__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_rs1[2]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_9__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[9]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_9__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_rs2[1]), .C2(Midori_rounds_sub_Sub_4_rs2[2]), 
        .A(Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_9__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_9__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_rs2[1]), .A2(Midori_rounds_sub_Sub_4_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_9__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_U3 ( .A(r[42]), 
        .B(r[43]), .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[2]), .B1(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[1]), .B2(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_10__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[11]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_4_rs2[1]), .C2(Midori_rounds_sub_Sub_4_rs2[2]), 
        .A(Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_4_rs2[1]), .A2(Midori_rounds_sub_Sub_4_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_rs1[3]), .B(Midori_rounds_sub_Sub_4_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_U1 ( .A(r[44]), 
        .B(r[43]), .Z(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_rs1[2]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[12]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_12__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_12__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_12__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_U3 ( .A(r[44]), 
        .B(r[45]), .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_4_rs2[5]), .B1(Midori_rounds_sub_Sub_4_rs2[4]), 
        .B2(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_13__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[14]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_rs1[3]), .B(Midori_rounds_sub_Sub_4_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_U1 ( .A(r[46]), 
        .B(r[45]), .Z(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_15__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_rs1[2]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_15__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[15]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_15__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_rs2[4]), .C2(Midori_rounds_sub_Sub_4_rs2[5]), 
        .A(Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_15__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_15__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_rs2[4]), .A2(Midori_rounds_sub_Sub_4_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_15__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[16]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_4_rs2[4]), .C2(Midori_rounds_sub_Sub_4_rs2[5]), 
        .A(Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_rs2[4]), .A2(Midori_rounds_sub_Sub_4_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_4_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_U1 ( .A(r[46]), 
        .B(r[47]), .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_16__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_U4 ( .A(r[42]), 
        .B(Midori_rounds_sub_Sub_4_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_n16) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_U3 ( .A(r[47]), 
        .B(Midori_rounds_sub_Sub_4_rs1[3]), .Z(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_n17) );
  AOI22_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_4_rs2[2]), .B1(Midori_rounds_sub_Sub_4_rs2[1]), 
        .B2(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_17__CF_Inst_n15) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_18__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_rs1[4]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_18__CF_Inst_n3), .Z(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_rs2[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_18__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_U2 ( .A(r[49]), 
        .B(r[48]), .Z(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_rs1[5]), .B(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_19__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_4_rs2[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_U4 ( .A(r[49]), 
        .B(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_U2 ( .A(r[50]), 
        .B(Midori_rounds_sub_Sub_4_rs2[0]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_rs1[4]), .B(Midori_rounds_sub_Sub_4_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_20__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_21__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_21__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_4_rs1[4]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[21]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_21__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_rs2[4]), .A2(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_U2 ( .A(r[51]), 
        .B(r[50]), .Z(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_rs1[5]), .B(Midori_rounds_sub_Sub_4_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_22__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[23]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_U4 ( .A(r[51]), 
        .B(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_U2 ( .A(r[52]), 
        .B(Midori_rounds_sub_Sub_4_S2_InAff_out3_reg[0]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_rs1[4]), .B(Midori_rounds_sub_Sub_4_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_23__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_24__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_24__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_4_rs1[4]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[24]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_rs2[4]), .A2(
        Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_24__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[25]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_rs2[4]), .A2(
        Midori_rounds_sub_Sub_4_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_U2 ( .A(r[53]), 
        .B(r[52]), .Z(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_rs1[5]), .B(Midori_rounds_sub_Sub_4_rs2[3]), 
        .ZN(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_4_rs2[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_U4 ( .A(r[53]), 
        .B(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_U2 ( .A(r[48]), 
        .B(Midori_rounds_sub_Sub_4_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_rs1[4]), .B(Midori_rounds_sub_Sub_4_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_4_S2_F_inst_Inst_26__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_1__Compression2_n2), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_1__Compression2_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_4_S2_F_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_4_S2_F_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result1[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_0__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_0__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[0]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_0__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_U2 ( .A(r[67]), 
        .B(r[66]), .Z(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_4_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_1__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_U2 ( .A(1'b0), .B(
        r[68]), .Z(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_U1 ( .A(1'b0), 
        .B(r[67]), .ZN(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_3__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_3__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_U2 ( .A(r[69]), 
        .B(r[68]), .Z(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_4_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_4__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[5]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_U2 ( .A(1'b0), .B(
        r[70]), .Z(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_U1 ( .A(1'b0), 
        .B(r[69]), .ZN(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_6__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_6__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[6]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_6__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_7__CF_Inst_U4 ( .A(1'b0), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_7__CF_Inst_n9), .Z(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_7__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_7__CF_Inst_n8), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_7__CF_Inst_n7), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_7__CF_Inst_n9) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_7__CF_Inst_n7) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_7__CF_Inst_U1 ( .A(r[70]), 
        .B(r[71]), .Z(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_7__CF_Inst_n8) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_U4 ( .A(r[71]), 
        .B(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_U2 ( .A(r[66]), 
        .B(Midori_rounds_sub_Sub_4_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_U1 ( .A(1'b0), .B(
        1'b0), .Z(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_8__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_9__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_9__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[9]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[1]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_U1 ( .A(r[54]), 
        .B(r[55]), .Z(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_10__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[11]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_U4 ( .A(r[55]), 
        .B(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_U2 ( .A(r[56]), 
        .B(Midori_rounds_sub_Sub_4_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_12__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[1]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_U1 ( .A(r[56]), 
        .B(r[57]), .Z(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_13__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[14]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_U4 ( .A(r[57]), 
        .B(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_U2 ( .A(r[58]), 
        .B(Midori_rounds_sub_Sub_4_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_15__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_15__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[15]) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_U2 ( .A(r[59]), 
        .B(r[58]), .Z(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_4_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_n13), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_n12), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_n12) );
  INV_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[1]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_U2 ( .A(r[59]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_n13)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_U1 ( .A(r[54]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_17__CF_Inst_n15)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_18__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_18__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[18]) );
  AOI21_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_18__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_18__CF_Inst_n6) );
  OAI21_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_18__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_U3 ( .A(r[60]), 
        .B(r[61]), .ZN(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[2]), .B1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[1]), .B2(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_19__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[20]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[1]), .C2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_U1 ( .A(r[62]), 
        .B(r[61]), .Z(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_20__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_21__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_21__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[21]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_21__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_21__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_U3 ( .A(r[62]), 
        .B(r[63]), .ZN(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[2]), .B1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[1]), .B2(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_22__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[23]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_U1 ( .A(r[64]), 
        .B(r[63]), .Z(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_23__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_24__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_24__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[24]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_24__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[25]) );
  OAI211_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[3]), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_n9), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_U1 ( .A(r[64]), 
        .B(r[65]), .ZN(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_25__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Out[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_U4 ( .A(r[60]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_n16)
         );
  XOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_U3 ( .A(r[65]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_n17)
         );
  AOI22_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[2]), .B1(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[18]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[18]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[18]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_4_S2_G_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_4_S2_G_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_InAff_out3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_S1_InAff_out3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_InAff_out3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_S1_InAff_out3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_InAff_out3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_S1_InAff_out3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_InAff_out3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_5_S1_InAff_out3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_S1_InAff_out2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_rs1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_S1_InAff_out2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_rs1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_S1_InAff_out2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_rs1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_5_S1_InAff_out2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_3_), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_S1_InAff_out1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_rs1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_S1_InAff_out1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_rs1[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_S1_InAff_out1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_rs1[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_5_S1_InAff_out1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_3_), .QN() );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_InputAffine_U3 ( .A(
        Midori_rounds_sub_Sub_5_S1_InAff_out3[1]), .B(Midori_rounds_n959), .Z(
        Midori_rounds_sub_Sub_5_S1_InAff_out3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_InputAffine_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_InAff_out2[1]), .B(Midori_rounds_n895), .Z(
        Midori_rounds_sub_Sub_5_S1_InAff_out2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_InputAffine_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_InAff_out1[1]), .B(Midori_rounds_n836), .Z(
        Midori_rounds_sub_Sub_5_S1_InAff_out1[3]) );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_rs1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_rs1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_0__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_rs2[0]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_0__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[0]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_0__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_rs1[1]), .C2(Midori_rounds_sub_Sub_5_rs1[2]), 
        .A(Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_0__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_0__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_rs1[1]), .A2(Midori_rounds_sub_Sub_5_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_0__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_5_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_U3 ( .A(r[0]), 
        .B(r[1]), .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_3_), .B2(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[1]), .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_1__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[2]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_5_rs1[1]), .C2(Midori_rounds_sub_Sub_5_rs1[2]), 
        .A(Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_5_rs1[1]), .A2(Midori_rounds_sub_Sub_5_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_rs2[1]), .B(Midori_rounds_sub_Sub_5_rs2[0]), 
        .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_U1 ( .A(r[2]), .B(
        r[1]), .Z(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_3__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_rs2[0]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_3__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[3]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_3__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_3__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_3__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_3__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_5_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_U3 ( .A(r[2]), 
        .B(r[3]), .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[3]), .B2(
        Midori_rounds_sub_Sub_5_rs1[4]), .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_5_rs1[5]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_4__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[5]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_rs2[1]), .B(Midori_rounds_sub_Sub_5_rs2[0]), 
        .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_U1 ( .A(r[4]), .B(
        r[3]), .Z(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_6__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_rs2[0]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_6__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[6]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_6__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_rs1[4]), .C2(Midori_rounds_sub_Sub_5_rs1[5]), 
        .A(Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_6__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_6__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_rs1[4]), .A2(Midori_rounds_sub_Sub_5_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_6__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[7]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_5_rs1[4]), .C2(Midori_rounds_sub_Sub_5_rs1[5]), 
        .A(Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_rs1[4]), .A2(Midori_rounds_sub_Sub_5_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_5_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_U1 ( .A(r[4]), 
        .B(r[5]), .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_7__CF_Inst_n9) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_n21), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_n20), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[8]) );
  OAI21_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_U5 ( .B1(
        Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_3_), .B2(
        Midori_rounds_sub_Sub_5_rs1[1]), .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_n19), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_n20) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_5_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_n19) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_n18), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_n17), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_n21) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_rs2[1]), .B(r[5]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_n17) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_rs2[0]), .B(r[0]), .Z(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_8__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_9__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_rs2[2]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_9__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[9]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_9__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_rs1[1]), .C2(Midori_rounds_sub_Sub_5_rs1[2]), 
        .A(Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_9__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_9__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_rs1[1]), .A2(Midori_rounds_sub_Sub_5_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_9__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_U3 ( .A(r[6]), 
        .B(r[7]), .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[2]), .B1(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_10__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[11]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_5_rs1[1]), .C2(Midori_rounds_sub_Sub_5_rs1[2]), 
        .A(Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_5_rs1[1]), .A2(Midori_rounds_sub_Sub_5_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_rs2[3]), .B(Midori_rounds_sub_Sub_5_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_U1 ( .A(r[8]), 
        .B(r[7]), .Z(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_rs2[2]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[12]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_12__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_12__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_12__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_U3 ( .A(r[8]), 
        .B(r[9]), .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_5_rs1[5]), .B1(Midori_rounds_sub_Sub_5_rs1[4]), 
        .B2(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_13__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[14]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_rs2[3]), .B(Midori_rounds_sub_Sub_5_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_U1 ( .A(r[10]), 
        .B(r[9]), .Z(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_15__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_rs2[2]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_15__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[15]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_15__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_rs1[4]), .C2(Midori_rounds_sub_Sub_5_rs1[5]), 
        .A(Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_15__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_15__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_rs1[4]), .A2(Midori_rounds_sub_Sub_5_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_15__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[16]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_5_rs1[4]), .C2(Midori_rounds_sub_Sub_5_rs1[5]), 
        .A(Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_rs1[4]), .A2(Midori_rounds_sub_Sub_5_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_5_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_U1 ( .A(r[10]), 
        .B(r[11]), .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_16__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_U4 ( .A(r[6]), 
        .B(Midori_rounds_sub_Sub_5_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_n16) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_U3 ( .A(r[11]), 
        .B(Midori_rounds_sub_Sub_5_rs2[3]), .Z(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_n17) );
  AOI22_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_5_rs1[2]), .B1(Midori_rounds_sub_Sub_5_rs1[1]), 
        .B2(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_17__CF_Inst_n15) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_18__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_rs2[4]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_18__CF_Inst_n3), .Z(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_rs1[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_18__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_U2 ( .A(r[13]), 
        .B(r[12]), .Z(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_rs2[5]), .B(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_19__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_5_rs1[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_U4 ( .A(r[13]), 
        .B(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_U2 ( .A(r[14]), 
        .B(Midori_rounds_sub_Sub_5_rs1[0]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_rs2[4]), .B(Midori_rounds_sub_Sub_5_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_20__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_21__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_21__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_5_rs2[4]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[21]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_21__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_rs1[4]), .A2(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_U2 ( .A(r[15]), 
        .B(r[14]), .Z(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_rs2[5]), .B(Midori_rounds_sub_Sub_5_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_22__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[23]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_U4 ( .A(r[15]), 
        .B(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_U2 ( .A(r[16]), 
        .B(Midori_rounds_sub_Sub_5_S1_InAff_out3_reg[0]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_rs2[4]), .B(Midori_rounds_sub_Sub_5_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_23__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_24__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_24__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_5_rs2[4]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[24]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_rs1[4]), .A2(
        Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_24__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[25]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_rs1[4]), .A2(
        Midori_rounds_sub_Sub_5_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_U2 ( .A(r[17]), 
        .B(r[16]), .Z(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_rs2[5]), .B(Midori_rounds_sub_Sub_5_rs1[3]), 
        .ZN(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_5_rs1[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_U4 ( .A(r[17]), 
        .B(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_U2 ( .A(r[12]), 
        .B(Midori_rounds_sub_Sub_5_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_rs2[4]), .B(Midori_rounds_sub_Sub_5_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_5_S1_F_inst_Inst_26__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_1__Compression2_n2), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_1__Compression2_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_5_S1_F_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_5_S1_F_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[53]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result1[53]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[53]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_0__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_0__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[0]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_0__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_U2 ( .A(r[31]), 
        .B(r[30]), .Z(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_5_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_1__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_U2 ( .A(1'b0), .B(
        r[32]), .Z(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_U1 ( .A(1'b0), 
        .B(r[31]), .ZN(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_3__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_3__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_U2 ( .A(r[33]), 
        .B(r[32]), .Z(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_5_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_4__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[5]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_U2 ( .A(1'b0), .B(
        r[34]), .Z(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_U1 ( .A(1'b0), 
        .B(r[33]), .ZN(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_6__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_6__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[6]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_6__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_7__CF_Inst_U4 ( .A(1'b0), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_7__CF_Inst_n9), .Z(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_7__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_7__CF_Inst_n8), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_7__CF_Inst_n7), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_7__CF_Inst_n9) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_7__CF_Inst_n7) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_7__CF_Inst_U1 ( .A(r[34]), 
        .B(r[35]), .Z(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_7__CF_Inst_n8) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_U4 ( .A(r[35]), 
        .B(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_U2 ( .A(r[30]), 
        .B(Midori_rounds_sub_Sub_5_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_U1 ( .A(1'b0), .B(
        1'b0), .Z(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_8__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_9__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_9__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[9]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[1]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_U1 ( .A(r[18]), 
        .B(r[19]), .Z(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_10__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[11]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_U4 ( .A(r[19]), 
        .B(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_U2 ( .A(r[20]), 
        .B(Midori_rounds_sub_Sub_5_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_12__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[1]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_U1 ( .A(r[20]), 
        .B(r[21]), .Z(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_13__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[14]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_U4 ( .A(r[21]), 
        .B(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_U2 ( .A(r[22]), 
        .B(Midori_rounds_sub_Sub_5_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_15__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_15__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[15]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_U2 ( .A(r[23]), 
        .B(r[22]), .Z(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_5_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_n13), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_n12), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_n12) );
  INV_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[1]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_U2 ( .A(r[23]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_n13)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_U1 ( .A(r[18]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_17__CF_Inst_n15)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_18__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_18__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[18]) );
  AOI21_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_18__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_18__CF_Inst_n6) );
  OAI21_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_18__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_U3 ( .A(r[24]), 
        .B(r[25]), .ZN(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[2]), .B1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[1]), .B2(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_19__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[20]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[1]), .C2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_U1 ( .A(r[26]), 
        .B(r[25]), .Z(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_20__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_21__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_21__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[21]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_21__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_21__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_U3 ( .A(r[26]), 
        .B(r[27]), .ZN(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[2]), .B1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[1]), .B2(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_22__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[23]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_U1 ( .A(r[28]), 
        .B(r[27]), .Z(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_23__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_24__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_24__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[24]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_24__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[25]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[3]), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_n9), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_U1 ( .A(r[28]), 
        .B(r[29]), .ZN(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_25__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Out[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_U4 ( .A(r[24]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_n16)
         );
  XOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_U3 ( .A(r[29]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_n17)
         );
  AOI22_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[2]), .B1(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[52]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[52]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[52]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[54]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[54]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[54]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[55]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[55]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[55]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_5_S1_G_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_5_S1_G_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_InAff_out3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_S2_InAff_out3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_InAff_out3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_S2_InAff_out3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_InAff_out3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_S2_InAff_out3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_InAff_out3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_5_S2_InAff_out3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_S2_InAff_out2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_rs2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_S2_InAff_out2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_rs2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_S2_InAff_out2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_rs2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_5_S2_InAff_out2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_3_), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_S2_InAff_out1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_rs2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_S2_InAff_out1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_rs2[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_S2_InAff_out1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_rs2[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_5_S2_InAff_out1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_3_), .QN() );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_InputAffine_U3 ( .A(
        Midori_rounds_sub_Sub_5_S2_InAff_out3[1]), .B(Midori_rounds_n963), .Z(
        Midori_rounds_sub_Sub_5_S2_InAff_out3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_InputAffine_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_InAff_out2[1]), .B(Midori_rounds_n899), .Z(
        Midori_rounds_sub_Sub_5_S2_InAff_out2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_InputAffine_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_InAff_out1[1]), .B(Midori_rounds_n839), .Z(
        Midori_rounds_sub_Sub_5_S2_InAff_out1[3]) );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_rs2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_rs2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_0__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_rs1[0]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_0__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[0]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_0__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_rs2[1]), .C2(Midori_rounds_sub_Sub_5_rs2[2]), 
        .A(Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_0__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_0__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_rs2[1]), .A2(Midori_rounds_sub_Sub_5_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_0__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_5_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_U3 ( .A(r[36]), 
        .B(r[37]), .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_3_), .B2(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[1]), .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_1__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[2]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_5_rs2[1]), .C2(Midori_rounds_sub_Sub_5_rs2[2]), 
        .A(Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_5_rs2[1]), .A2(Midori_rounds_sub_Sub_5_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_rs1[1]), .B(Midori_rounds_sub_Sub_5_rs1[0]), 
        .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_U1 ( .A(r[38]), 
        .B(r[37]), .Z(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_3__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_rs1[0]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_3__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[3]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_3__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_3__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_3__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_3__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_5_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_U3 ( .A(r[38]), 
        .B(r[39]), .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[3]), .B2(
        Midori_rounds_sub_Sub_5_rs2[4]), .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_5_rs2[5]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_4__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[5]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_rs1[1]), .B(Midori_rounds_sub_Sub_5_rs1[0]), 
        .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_U1 ( .A(r[40]), 
        .B(r[39]), .Z(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_6__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_rs1[0]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_6__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[6]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_6__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_rs2[4]), .C2(Midori_rounds_sub_Sub_5_rs2[5]), 
        .A(Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_6__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_6__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_rs2[4]), .A2(Midori_rounds_sub_Sub_5_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_6__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[7]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_5_rs2[4]), .C2(Midori_rounds_sub_Sub_5_rs2[5]), 
        .A(Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_rs2[4]), .A2(Midori_rounds_sub_Sub_5_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_5_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_U1 ( .A(r[40]), 
        .B(r[41]), .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_7__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_n21), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_n20), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[8]) );
  OAI21_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_U5 ( .B1(
        Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_3_), .B2(
        Midori_rounds_sub_Sub_5_rs2[1]), .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_n19), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_n20) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_5_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_n19) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_n18), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_n17), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_n21) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_rs1[1]), .B(r[41]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_n17) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_rs1[0]), .B(r[36]), .Z(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_8__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_9__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_rs1[2]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_9__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[9]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_9__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_rs2[1]), .C2(Midori_rounds_sub_Sub_5_rs2[2]), 
        .A(Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_9__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_9__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_rs2[1]), .A2(Midori_rounds_sub_Sub_5_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_9__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_U3 ( .A(r[42]), 
        .B(r[43]), .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[2]), .B1(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[1]), .B2(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_10__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[11]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_5_rs2[1]), .C2(Midori_rounds_sub_Sub_5_rs2[2]), 
        .A(Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_5_rs2[1]), .A2(Midori_rounds_sub_Sub_5_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_rs1[3]), .B(Midori_rounds_sub_Sub_5_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_U1 ( .A(r[44]), 
        .B(r[43]), .Z(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_rs1[2]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[12]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_12__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_12__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_12__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_U3 ( .A(r[44]), 
        .B(r[45]), .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_5_rs2[5]), .B1(Midori_rounds_sub_Sub_5_rs2[4]), 
        .B2(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_13__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[14]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_rs1[3]), .B(Midori_rounds_sub_Sub_5_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_U1 ( .A(r[46]), 
        .B(r[45]), .Z(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_15__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_rs1[2]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_15__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[15]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_15__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_rs2[4]), .C2(Midori_rounds_sub_Sub_5_rs2[5]), 
        .A(Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_15__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_15__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_rs2[4]), .A2(Midori_rounds_sub_Sub_5_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_15__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[16]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_5_rs2[4]), .C2(Midori_rounds_sub_Sub_5_rs2[5]), 
        .A(Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_rs2[4]), .A2(Midori_rounds_sub_Sub_5_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_5_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_U1 ( .A(r[46]), 
        .B(r[47]), .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_16__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_U4 ( .A(r[42]), 
        .B(Midori_rounds_sub_Sub_5_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_n16) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_U3 ( .A(r[47]), 
        .B(Midori_rounds_sub_Sub_5_rs1[3]), .Z(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_n17) );
  AOI22_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_5_rs2[2]), .B1(Midori_rounds_sub_Sub_5_rs2[1]), 
        .B2(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_17__CF_Inst_n15) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_18__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_rs1[4]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_18__CF_Inst_n3), .Z(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_rs2[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_18__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_U2 ( .A(r[49]), 
        .B(r[48]), .Z(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_rs1[5]), .B(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_19__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_5_rs2[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_U4 ( .A(r[49]), 
        .B(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_U2 ( .A(r[50]), 
        .B(Midori_rounds_sub_Sub_5_rs2[0]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_rs1[4]), .B(Midori_rounds_sub_Sub_5_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_20__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_21__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_21__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_5_rs1[4]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[21]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_21__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_rs2[4]), .A2(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_U2 ( .A(r[51]), 
        .B(r[50]), .Z(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_rs1[5]), .B(Midori_rounds_sub_Sub_5_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_22__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[23]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_U4 ( .A(r[51]), 
        .B(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_U2 ( .A(r[52]), 
        .B(Midori_rounds_sub_Sub_5_S2_InAff_out3_reg[0]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_rs1[4]), .B(Midori_rounds_sub_Sub_5_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_23__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_24__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_24__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_5_rs1[4]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[24]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_rs2[4]), .A2(
        Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_24__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[25]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_rs2[4]), .A2(
        Midori_rounds_sub_Sub_5_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_U2 ( .A(r[53]), 
        .B(r[52]), .Z(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_rs1[5]), .B(Midori_rounds_sub_Sub_5_rs2[3]), 
        .ZN(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_5_rs2[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_U4 ( .A(r[53]), 
        .B(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_U2 ( .A(r[48]), 
        .B(Midori_rounds_sub_Sub_5_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_rs1[4]), .B(Midori_rounds_sub_Sub_5_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_5_S2_F_inst_Inst_26__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_1__Compression2_n2), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_1__Compression2_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_5_S2_F_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_5_S2_F_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[41]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result1[41]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[41]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_0__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_0__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[0]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_0__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_U2 ( .A(r[67]), 
        .B(r[66]), .Z(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_5_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_1__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_U2 ( .A(1'b0), .B(
        r[68]), .Z(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_U1 ( .A(1'b0), 
        .B(r[67]), .ZN(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_3__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_3__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_U2 ( .A(r[69]), 
        .B(r[68]), .Z(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_5_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_4__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[5]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_U2 ( .A(1'b0), .B(
        r[70]), .Z(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_U1 ( .A(1'b0), 
        .B(r[69]), .ZN(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_6__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_6__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[6]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_6__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_7__CF_Inst_U4 ( .A(1'b0), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_7__CF_Inst_n9), .Z(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_7__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_7__CF_Inst_n8), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_7__CF_Inst_n7), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_7__CF_Inst_n9) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_7__CF_Inst_n7) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_7__CF_Inst_U1 ( .A(r[70]), 
        .B(r[71]), .Z(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_7__CF_Inst_n8) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_U4 ( .A(r[71]), 
        .B(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_U2 ( .A(r[66]), 
        .B(Midori_rounds_sub_Sub_5_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_U1 ( .A(1'b0), .B(
        1'b0), .Z(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_8__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_9__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_9__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[9]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[1]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_U1 ( .A(r[54]), 
        .B(r[55]), .Z(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_10__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[11]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_U4 ( .A(r[55]), 
        .B(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_U2 ( .A(r[56]), 
        .B(Midori_rounds_sub_Sub_5_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_12__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[1]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_U1 ( .A(r[56]), 
        .B(r[57]), .Z(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_13__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[14]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_U4 ( .A(r[57]), 
        .B(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_U2 ( .A(r[58]), 
        .B(Midori_rounds_sub_Sub_5_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_15__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_15__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[15]) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_U2 ( .A(r[59]), 
        .B(r[58]), .Z(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_5_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_n13), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_n12), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_n12) );
  INV_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[1]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_U2 ( .A(r[59]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_n13)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_U1 ( .A(r[54]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_17__CF_Inst_n15)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_18__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_18__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[18]) );
  AOI21_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_18__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_18__CF_Inst_n6) );
  OAI21_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_18__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_U3 ( .A(r[60]), 
        .B(r[61]), .ZN(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[2]), .B1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[1]), .B2(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_19__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[20]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[1]), .C2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_U1 ( .A(r[62]), 
        .B(r[61]), .Z(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_20__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_21__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_21__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[21]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_21__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_21__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_U3 ( .A(r[62]), 
        .B(r[63]), .ZN(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[2]), .B1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[1]), .B2(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_22__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[23]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_U1 ( .A(r[64]), 
        .B(r[63]), .Z(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_23__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_24__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_24__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[24]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_24__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[25]) );
  OAI211_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[3]), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_n9), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_U1 ( .A(r[64]), 
        .B(r[65]), .ZN(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_25__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Out[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_U4 ( .A(r[60]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_n16)
         );
  XOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_U3 ( .A(r[65]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_n17)
         );
  AOI22_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[2]), .B1(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[40]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[40]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[40]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[42]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[42]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[42]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[43]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[43]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[43]) );
  XNOR2_X1 Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_5_S2_G_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_5_S2_G_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_InAff_out3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_S1_InAff_out3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_InAff_out3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_S1_InAff_out3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_InAff_out3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_S1_InAff_out3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_InAff_out3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_6_S1_InAff_out3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_S1_InAff_out2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_rs1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_S1_InAff_out2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_rs1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_S1_InAff_out2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_rs1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_6_S1_InAff_out2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_3_), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_S1_InAff_out1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_rs1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_S1_InAff_out1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_rs1[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_S1_InAff_out1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_rs1[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_6_S1_InAff_out1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_3_), .QN() );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_InputAffine_U3 ( .A(
        Midori_rounds_sub_Sub_6_S1_InAff_out3[1]), .B(Midori_rounds_n967), .Z(
        Midori_rounds_sub_Sub_6_S1_InAff_out3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_InputAffine_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_InAff_out2[1]), .B(Midori_rounds_n903), .Z(
        Midori_rounds_sub_Sub_6_S1_InAff_out2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_InputAffine_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_InAff_out1[1]), .B(Midori_rounds_n842), .Z(
        Midori_rounds_sub_Sub_6_S1_InAff_out1[3]) );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_rs1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_rs1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_0__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_rs2[0]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_0__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[0]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_0__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_rs1[1]), .C2(Midori_rounds_sub_Sub_6_rs1[2]), 
        .A(Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_0__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_0__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_rs1[1]), .A2(Midori_rounds_sub_Sub_6_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_0__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_6_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_U3 ( .A(r[0]), 
        .B(r[1]), .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_3_), .B2(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[1]), .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_1__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[2]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_6_rs1[1]), .C2(Midori_rounds_sub_Sub_6_rs1[2]), 
        .A(Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_6_rs1[1]), .A2(Midori_rounds_sub_Sub_6_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_rs2[1]), .B(Midori_rounds_sub_Sub_6_rs2[0]), 
        .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_U1 ( .A(r[2]), .B(
        r[1]), .Z(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_3__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_rs2[0]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_3__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[3]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_3__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_3__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_3__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_3__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_6_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_U3 ( .A(r[2]), 
        .B(r[3]), .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[3]), .B2(
        Midori_rounds_sub_Sub_6_rs1[4]), .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_6_rs1[5]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_4__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[5]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_rs2[1]), .B(Midori_rounds_sub_Sub_6_rs2[0]), 
        .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_U1 ( .A(r[4]), .B(
        r[3]), .Z(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_6__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_rs2[0]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_6__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[6]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_6__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_rs1[4]), .C2(Midori_rounds_sub_Sub_6_rs1[5]), 
        .A(Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_6__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_6__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_rs1[4]), .A2(Midori_rounds_sub_Sub_6_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_6__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[7]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_6_rs1[4]), .C2(Midori_rounds_sub_Sub_6_rs1[5]), 
        .A(Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_rs1[4]), .A2(Midori_rounds_sub_Sub_6_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_6_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_U1 ( .A(r[4]), 
        .B(r[5]), .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_7__CF_Inst_n9) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_n21), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_n20), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[8]) );
  OAI21_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_U5 ( .B1(
        Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_3_), .B2(
        Midori_rounds_sub_Sub_6_rs1[1]), .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_n19), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_n20) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_6_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_n19) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_n18), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_n17), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_n21) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_rs2[1]), .B(r[5]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_n17) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_rs2[0]), .B(r[0]), .Z(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_8__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_9__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_rs2[2]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_9__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[9]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_9__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_rs1[1]), .C2(Midori_rounds_sub_Sub_6_rs1[2]), 
        .A(Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_9__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_9__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_rs1[1]), .A2(Midori_rounds_sub_Sub_6_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_9__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_U3 ( .A(r[6]), 
        .B(r[7]), .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[2]), .B1(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_10__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[11]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_6_rs1[1]), .C2(Midori_rounds_sub_Sub_6_rs1[2]), 
        .A(Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_6_rs1[1]), .A2(Midori_rounds_sub_Sub_6_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_rs2[3]), .B(Midori_rounds_sub_Sub_6_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_U1 ( .A(r[8]), 
        .B(r[7]), .Z(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_rs2[2]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[12]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_12__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_12__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_12__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_U3 ( .A(r[8]), 
        .B(r[9]), .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_6_rs1[5]), .B1(Midori_rounds_sub_Sub_6_rs1[4]), 
        .B2(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_13__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[14]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_rs2[3]), .B(Midori_rounds_sub_Sub_6_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_U1 ( .A(r[10]), 
        .B(r[9]), .Z(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_15__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_rs2[2]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_15__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[15]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_15__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_rs1[4]), .C2(Midori_rounds_sub_Sub_6_rs1[5]), 
        .A(Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_15__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_15__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_rs1[4]), .A2(Midori_rounds_sub_Sub_6_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_15__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[16]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_6_rs1[4]), .C2(Midori_rounds_sub_Sub_6_rs1[5]), 
        .A(Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_rs1[4]), .A2(Midori_rounds_sub_Sub_6_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_6_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_U1 ( .A(r[10]), 
        .B(r[11]), .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_16__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_U4 ( .A(r[6]), 
        .B(Midori_rounds_sub_Sub_6_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_n16) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_U3 ( .A(r[11]), 
        .B(Midori_rounds_sub_Sub_6_rs2[3]), .Z(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_n17) );
  AOI22_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_6_rs1[2]), .B1(Midori_rounds_sub_Sub_6_rs1[1]), 
        .B2(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_17__CF_Inst_n15) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_18__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_rs2[4]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_18__CF_Inst_n3), .Z(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_rs1[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_18__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_U2 ( .A(r[13]), 
        .B(r[12]), .Z(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_rs2[5]), .B(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_19__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_6_rs1[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_U4 ( .A(r[13]), 
        .B(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_U2 ( .A(r[14]), 
        .B(Midori_rounds_sub_Sub_6_rs1[0]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_rs2[4]), .B(Midori_rounds_sub_Sub_6_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_20__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_21__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_21__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_6_rs2[4]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[21]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_21__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_rs1[4]), .A2(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_U2 ( .A(r[15]), 
        .B(r[14]), .Z(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_rs2[5]), .B(Midori_rounds_sub_Sub_6_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_22__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[23]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_U4 ( .A(r[15]), 
        .B(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_U2 ( .A(r[16]), 
        .B(Midori_rounds_sub_Sub_6_S1_InAff_out3_reg[0]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_rs2[4]), .B(Midori_rounds_sub_Sub_6_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_23__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_24__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_24__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_6_rs2[4]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[24]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_rs1[4]), .A2(
        Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_24__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[25]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_rs1[4]), .A2(
        Midori_rounds_sub_Sub_6_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_U2 ( .A(r[17]), 
        .B(r[16]), .Z(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_rs2[5]), .B(Midori_rounds_sub_Sub_6_rs1[3]), 
        .ZN(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_6_rs1[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_U4 ( .A(r[17]), 
        .B(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_U2 ( .A(r[12]), 
        .B(Midori_rounds_sub_Sub_6_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_rs2[4]), .B(Midori_rounds_sub_Sub_6_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_6_S1_F_inst_Inst_26__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_1__Compression2_n2), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_1__Compression2_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_6_S1_F_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_6_S1_F_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result1[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_0__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_0__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[0]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_0__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_U2 ( .A(r[31]), 
        .B(r[30]), .Z(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_6_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_1__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_U2 ( .A(1'b0), .B(
        r[32]), .Z(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_U1 ( .A(1'b0), 
        .B(r[31]), .ZN(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_3__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_3__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_U2 ( .A(r[33]), 
        .B(r[32]), .Z(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_6_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_4__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[5]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_U2 ( .A(1'b0), .B(
        r[34]), .Z(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_U1 ( .A(1'b0), 
        .B(r[33]), .ZN(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_6__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_6__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[6]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_6__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_7__CF_Inst_U4 ( .A(1'b0), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_7__CF_Inst_n9), .Z(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_7__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_7__CF_Inst_n8), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_7__CF_Inst_n7), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_7__CF_Inst_n9) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_7__CF_Inst_n7) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_7__CF_Inst_U1 ( .A(r[34]), 
        .B(r[35]), .Z(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_7__CF_Inst_n8) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_U4 ( .A(r[35]), 
        .B(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_U2 ( .A(r[30]), 
        .B(Midori_rounds_sub_Sub_6_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_U1 ( .A(1'b0), .B(
        1'b0), .Z(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_8__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_9__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_9__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[9]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[1]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_U1 ( .A(r[18]), 
        .B(r[19]), .Z(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_10__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[11]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_U4 ( .A(r[19]), 
        .B(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_U2 ( .A(r[20]), 
        .B(Midori_rounds_sub_Sub_6_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_12__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[1]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_U1 ( .A(r[20]), 
        .B(r[21]), .Z(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_13__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[14]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_U4 ( .A(r[21]), 
        .B(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_U2 ( .A(r[22]), 
        .B(Midori_rounds_sub_Sub_6_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_15__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_15__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[15]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_U2 ( .A(r[23]), 
        .B(r[22]), .Z(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_6_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_n13), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_n12), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_n12) );
  INV_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[1]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_U2 ( .A(r[23]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_n13)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_U1 ( .A(r[18]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_17__CF_Inst_n15)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_18__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_18__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[18]) );
  AOI21_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_18__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_18__CF_Inst_n6) );
  OAI21_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_18__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_U3 ( .A(r[24]), 
        .B(r[25]), .ZN(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[2]), .B1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[1]), .B2(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_19__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[20]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[1]), .C2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_U1 ( .A(r[26]), 
        .B(r[25]), .Z(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_20__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_21__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_21__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[21]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_21__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_21__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_U3 ( .A(r[26]), 
        .B(r[27]), .ZN(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[2]), .B1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[1]), .B2(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_22__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[23]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_U1 ( .A(r[28]), 
        .B(r[27]), .Z(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_23__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_24__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_24__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[24]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_24__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[25]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[3]), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_n9), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_U1 ( .A(r[28]), 
        .B(r[29]), .ZN(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_25__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Out[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_U4 ( .A(r[24]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_n16)
         );
  XOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_U3 ( .A(r[29]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_n17)
         );
  AOI22_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[2]), .B1(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[24]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[24]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[24]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[27]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[27]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[27]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_6_S1_G_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_6_S1_G_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_InAff_out3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_S2_InAff_out3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_InAff_out3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_S2_InAff_out3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_InAff_out3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_S2_InAff_out3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_InAff_out3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_6_S2_InAff_out3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_S2_InAff_out2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_rs2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_S2_InAff_out2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_rs2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_S2_InAff_out2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_rs2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_6_S2_InAff_out2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_3_), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_S2_InAff_out1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_rs2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_S2_InAff_out1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_rs2[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_S2_InAff_out1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_rs2[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_6_S2_InAff_out1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_3_), .QN() );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_InputAffine_U3 ( .A(
        Midori_rounds_sub_Sub_6_S2_InAff_out3[1]), .B(Midori_rounds_n971), .Z(
        Midori_rounds_sub_Sub_6_S2_InAff_out3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_InputAffine_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_InAff_out2[1]), .B(Midori_rounds_n907), .Z(
        Midori_rounds_sub_Sub_6_S2_InAff_out2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_InputAffine_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_InAff_out1[1]), .B(Midori_rounds_n845), .Z(
        Midori_rounds_sub_Sub_6_S2_InAff_out1[3]) );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_rs2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_rs2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_0__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_rs1[0]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_0__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[0]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_0__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_rs2[1]), .C2(Midori_rounds_sub_Sub_6_rs2[2]), 
        .A(Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_0__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_0__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_rs2[1]), .A2(Midori_rounds_sub_Sub_6_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_0__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_6_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_U3 ( .A(r[36]), 
        .B(r[37]), .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_3_), .B2(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[1]), .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_1__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[2]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_6_rs2[1]), .C2(Midori_rounds_sub_Sub_6_rs2[2]), 
        .A(Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_6_rs2[1]), .A2(Midori_rounds_sub_Sub_6_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_rs1[1]), .B(Midori_rounds_sub_Sub_6_rs1[0]), 
        .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_U1 ( .A(r[38]), 
        .B(r[37]), .Z(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_3__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_rs1[0]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_3__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[3]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_3__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_3__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_3__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_3__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_6_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_U3 ( .A(r[38]), 
        .B(r[39]), .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[3]), .B2(
        Midori_rounds_sub_Sub_6_rs2[4]), .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_6_rs2[5]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_4__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[5]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_rs1[1]), .B(Midori_rounds_sub_Sub_6_rs1[0]), 
        .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_U1 ( .A(r[40]), 
        .B(r[39]), .Z(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_6__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_rs1[0]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_6__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[6]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_6__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_rs2[4]), .C2(Midori_rounds_sub_Sub_6_rs2[5]), 
        .A(Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_6__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_6__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_rs2[4]), .A2(Midori_rounds_sub_Sub_6_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_6__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[7]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_6_rs2[4]), .C2(Midori_rounds_sub_Sub_6_rs2[5]), 
        .A(Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_rs2[4]), .A2(Midori_rounds_sub_Sub_6_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_6_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_U1 ( .A(r[40]), 
        .B(r[41]), .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_7__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_n21), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_n20), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[8]) );
  OAI21_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_U5 ( .B1(
        Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_3_), .B2(
        Midori_rounds_sub_Sub_6_rs2[1]), .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_n19), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_n20) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_6_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_n19) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_n18), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_n17), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_n21) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_rs1[1]), .B(r[41]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_n17) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_rs1[0]), .B(r[36]), .Z(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_8__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_9__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_rs1[2]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_9__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[9]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_9__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_rs2[1]), .C2(Midori_rounds_sub_Sub_6_rs2[2]), 
        .A(Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_9__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_9__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_rs2[1]), .A2(Midori_rounds_sub_Sub_6_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_9__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_U3 ( .A(r[42]), 
        .B(r[43]), .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[2]), .B1(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[1]), .B2(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_10__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[11]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_6_rs2[1]), .C2(Midori_rounds_sub_Sub_6_rs2[2]), 
        .A(Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_6_rs2[1]), .A2(Midori_rounds_sub_Sub_6_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_rs1[3]), .B(Midori_rounds_sub_Sub_6_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_U1 ( .A(r[44]), 
        .B(r[43]), .Z(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_rs1[2]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[12]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_12__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_12__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_12__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_U3 ( .A(r[44]), 
        .B(r[45]), .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_6_rs2[5]), .B1(Midori_rounds_sub_Sub_6_rs2[4]), 
        .B2(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_13__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[14]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_rs1[3]), .B(Midori_rounds_sub_Sub_6_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_U1 ( .A(r[46]), 
        .B(r[45]), .Z(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_15__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_rs1[2]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_15__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[15]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_15__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_rs2[4]), .C2(Midori_rounds_sub_Sub_6_rs2[5]), 
        .A(Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_15__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_15__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_rs2[4]), .A2(Midori_rounds_sub_Sub_6_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_15__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[16]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_6_rs2[4]), .C2(Midori_rounds_sub_Sub_6_rs2[5]), 
        .A(Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_rs2[4]), .A2(Midori_rounds_sub_Sub_6_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_6_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_U1 ( .A(r[46]), 
        .B(r[47]), .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_16__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_U4 ( .A(r[42]), 
        .B(Midori_rounds_sub_Sub_6_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_n16) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_U3 ( .A(r[47]), 
        .B(Midori_rounds_sub_Sub_6_rs1[3]), .Z(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_n17) );
  AOI22_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_6_rs2[2]), .B1(Midori_rounds_sub_Sub_6_rs2[1]), 
        .B2(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_17__CF_Inst_n15) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_18__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_rs1[4]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_18__CF_Inst_n3), .Z(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_rs2[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_18__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_U2 ( .A(r[49]), 
        .B(r[48]), .Z(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_rs1[5]), .B(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_19__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_6_rs2[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_U4 ( .A(r[49]), 
        .B(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_U2 ( .A(r[50]), 
        .B(Midori_rounds_sub_Sub_6_rs2[0]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_rs1[4]), .B(Midori_rounds_sub_Sub_6_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_20__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_21__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_21__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_6_rs1[4]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[21]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_21__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_rs2[4]), .A2(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_U2 ( .A(r[51]), 
        .B(r[50]), .Z(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_rs1[5]), .B(Midori_rounds_sub_Sub_6_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_22__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[23]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_U4 ( .A(r[51]), 
        .B(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_U2 ( .A(r[52]), 
        .B(Midori_rounds_sub_Sub_6_S2_InAff_out3_reg[0]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_rs1[4]), .B(Midori_rounds_sub_Sub_6_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_23__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_24__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_24__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_6_rs1[4]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[24]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_rs2[4]), .A2(
        Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_24__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[25]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_rs2[4]), .A2(
        Midori_rounds_sub_Sub_6_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_U2 ( .A(r[53]), 
        .B(r[52]), .Z(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_rs1[5]), .B(Midori_rounds_sub_Sub_6_rs2[3]), 
        .ZN(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_6_rs2[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_U4 ( .A(r[53]), 
        .B(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_U2 ( .A(r[48]), 
        .B(Midori_rounds_sub_Sub_6_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_rs1[4]), .B(Midori_rounds_sub_Sub_6_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_6_S2_F_inst_Inst_26__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_1__Compression2_n2), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_1__Compression2_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_6_S2_F_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_6_S2_F_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result1[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_0__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_0__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[0]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_0__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_U2 ( .A(r[67]), 
        .B(r[66]), .Z(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_6_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_1__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_U2 ( .A(1'b0), .B(
        r[68]), .Z(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_U1 ( .A(1'b0), 
        .B(r[67]), .ZN(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_3__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_3__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_U2 ( .A(r[69]), 
        .B(r[68]), .Z(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_6_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_4__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[5]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_U2 ( .A(1'b0), .B(
        r[70]), .Z(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_U1 ( .A(1'b0), 
        .B(r[69]), .ZN(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_6__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_6__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[6]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_6__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_7__CF_Inst_U4 ( .A(1'b0), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_7__CF_Inst_n9), .Z(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_7__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_7__CF_Inst_n8), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_7__CF_Inst_n7), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_7__CF_Inst_n9) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_7__CF_Inst_n7) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_7__CF_Inst_U1 ( .A(r[70]), 
        .B(r[71]), .Z(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_7__CF_Inst_n8) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_U4 ( .A(r[71]), 
        .B(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_U2 ( .A(r[66]), 
        .B(Midori_rounds_sub_Sub_6_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_U1 ( .A(1'b0), .B(
        1'b0), .Z(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_8__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_9__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_9__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[9]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[1]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_U1 ( .A(r[54]), 
        .B(r[55]), .Z(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_10__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[11]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_U4 ( .A(r[55]), 
        .B(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_U2 ( .A(r[56]), 
        .B(Midori_rounds_sub_Sub_6_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_12__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[1]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_U1 ( .A(r[56]), 
        .B(r[57]), .Z(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_13__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[14]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_U4 ( .A(r[57]), 
        .B(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_U2 ( .A(r[58]), 
        .B(Midori_rounds_sub_Sub_6_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_15__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_15__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[15]) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_U2 ( .A(r[59]), 
        .B(r[58]), .Z(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_6_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_n13), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_n12), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_n12) );
  INV_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[1]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_U2 ( .A(r[59]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_n13)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_U1 ( .A(r[54]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_17__CF_Inst_n15)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_18__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_18__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[18]) );
  AOI21_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_18__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_18__CF_Inst_n6) );
  OAI21_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_18__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_U3 ( .A(r[60]), 
        .B(r[61]), .ZN(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[2]), .B1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[1]), .B2(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_19__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[20]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[1]), .C2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_U1 ( .A(r[62]), 
        .B(r[61]), .Z(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_20__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_21__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_21__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[21]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_21__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_21__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_U3 ( .A(r[62]), 
        .B(r[63]), .ZN(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[2]), .B1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[1]), .B2(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_22__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[23]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_U1 ( .A(r[64]), 
        .B(r[63]), .Z(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_23__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_24__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_24__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[24]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_24__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[25]) );
  OAI211_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[3]), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_n9), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_U1 ( .A(r[64]), 
        .B(r[65]), .ZN(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_25__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Out[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_U4 ( .A(r[60]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_n16)
         );
  XOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_U3 ( .A(r[65]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_n17)
         );
  AOI22_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[2]), .B1(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[6]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[6]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[6]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_6_S2_G_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_6_S2_G_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_InAff_out3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_S1_InAff_out3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_InAff_out3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_S1_InAff_out3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_InAff_out3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_S1_InAff_out3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_InAff_out3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_7_S1_InAff_out3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_S1_InAff_out2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_rs1[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_S1_InAff_out2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_rs1[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_S1_InAff_out2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_rs1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_7_S1_InAff_out2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_3_), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_S1_InAff_out1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_rs1[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_S1_InAff_out1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_rs1[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_S1_InAff_out1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_rs1[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_7_S1_InAff_out1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_3_), .QN() );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_InputAffine_U3 ( .A(
        Midori_rounds_sub_Sub_7_S1_InAff_out3[1]), .B(Midori_rounds_n975), .Z(
        Midori_rounds_sub_Sub_7_S1_InAff_out3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_InputAffine_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_InAff_out2[1]), .B(Midori_rounds_n911), .Z(
        Midori_rounds_sub_Sub_7_S1_InAff_out2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_InputAffine_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_InAff_out1[1]), .B(Midori_rounds_n848), .Z(
        Midori_rounds_sub_Sub_7_S1_InAff_out1[3]) );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_rs1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_rs1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_0__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_rs2[0]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_0__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[0]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_0__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_rs1[1]), .C2(Midori_rounds_sub_Sub_7_rs1[2]), 
        .A(Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_0__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_0__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_rs1[1]), .A2(Midori_rounds_sub_Sub_7_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_0__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_7_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_U3 ( .A(r[0]), 
        .B(r[1]), .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_3_), .B2(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[1]), .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_1__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[2]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_7_rs1[1]), .C2(Midori_rounds_sub_Sub_7_rs1[2]), 
        .A(Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_7_rs1[1]), .A2(Midori_rounds_sub_Sub_7_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_rs2[1]), .B(Midori_rounds_sub_Sub_7_rs2[0]), 
        .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_U1 ( .A(r[2]), .B(
        r[1]), .Z(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_2__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_3__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_rs2[0]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_3__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[3]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_3__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_3__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_3__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_3__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_7_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_U3 ( .A(r[2]), 
        .B(r[3]), .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[3]), .B2(
        Midori_rounds_sub_Sub_7_rs1[4]), .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_7_rs1[5]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_4__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[5]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_rs2[1]), .B(Midori_rounds_sub_Sub_7_rs2[0]), 
        .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_U1 ( .A(r[4]), .B(
        r[3]), .Z(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_5__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_6__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_rs2[0]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_6__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[6]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_6__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_rs1[4]), .C2(Midori_rounds_sub_Sub_7_rs1[5]), 
        .A(Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_6__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_6__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_rs1[4]), .A2(Midori_rounds_sub_Sub_7_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_6__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[7]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_7_rs1[4]), .C2(Midori_rounds_sub_Sub_7_rs1[5]), 
        .A(Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_rs1[4]), .A2(Midori_rounds_sub_Sub_7_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_7_rs2[1]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_U1 ( .A(r[4]), 
        .B(r[5]), .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_7__CF_Inst_n9) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_n21), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_n20), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[8]) );
  OAI21_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_U5 ( .B1(
        Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_3_), .B2(
        Midori_rounds_sub_Sub_7_rs1[1]), .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_n19), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_n20) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_7_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_n19) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_n18), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_n17), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_n21) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_rs2[1]), .B(r[5]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_n17) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_rs2[0]), .B(r[0]), .Z(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_8__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_9__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_rs2[2]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_9__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[9]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_9__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_rs1[1]), .C2(Midori_rounds_sub_Sub_7_rs1[2]), 
        .A(Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_9__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_9__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_rs1[1]), .A2(Midori_rounds_sub_Sub_7_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_9__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_U3 ( .A(r[6]), 
        .B(r[7]), .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[2]), .B1(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_10__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[11]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_7_rs1[1]), .C2(Midori_rounds_sub_Sub_7_rs1[2]), 
        .A(Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_7_rs1[1]), .A2(Midori_rounds_sub_Sub_7_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_rs2[3]), .B(Midori_rounds_sub_Sub_7_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_U1 ( .A(r[8]), 
        .B(r[7]), .Z(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_rs2[2]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[12]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_12__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_12__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_12__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_U3 ( .A(r[8]), 
        .B(r[9]), .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_7_rs1[5]), .B1(Midori_rounds_sub_Sub_7_rs1[4]), 
        .B2(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_13__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[14]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_rs2[3]), .B(Midori_rounds_sub_Sub_7_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_U1 ( .A(r[10]), 
        .B(r[9]), .Z(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_15__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_rs2[2]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_15__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[15]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_15__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_rs1[4]), .C2(Midori_rounds_sub_Sub_7_rs1[5]), 
        .A(Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_15__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_15__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_rs1[4]), .A2(Midori_rounds_sub_Sub_7_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_15__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[16]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_7_rs1[4]), .C2(Midori_rounds_sub_Sub_7_rs1[5]), 
        .A(Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_rs1[4]), .A2(Midori_rounds_sub_Sub_7_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_7_rs2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_U1 ( .A(r[10]), 
        .B(r[11]), .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_16__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_U4 ( .A(r[6]), 
        .B(Midori_rounds_sub_Sub_7_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_n16) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_U3 ( .A(r[11]), 
        .B(Midori_rounds_sub_Sub_7_rs2[3]), .Z(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_n17) );
  AOI22_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_7_rs1[2]), .B1(Midori_rounds_sub_Sub_7_rs1[1]), 
        .B2(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_17__CF_Inst_n15) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_18__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_rs2[4]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_18__CF_Inst_n3), .Z(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_rs1[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_18__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_U2 ( .A(r[13]), 
        .B(r[12]), .Z(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_rs2[5]), .B(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_19__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_7_rs1[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_U4 ( .A(r[13]), 
        .B(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_U2 ( .A(r[14]), 
        .B(Midori_rounds_sub_Sub_7_rs1[0]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_rs2[4]), .B(Midori_rounds_sub_Sub_7_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_20__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_21__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_21__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_7_rs2[4]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[21]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_21__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_rs1[4]), .A2(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_U2 ( .A(r[15]), 
        .B(r[14]), .Z(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_rs2[5]), .B(Midori_rounds_sub_Sub_7_rs1[5]), 
        .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_22__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[23]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_U4 ( .A(r[15]), 
        .B(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_U2 ( .A(r[16]), 
        .B(Midori_rounds_sub_Sub_7_S1_InAff_out3_reg[0]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_rs2[4]), .B(Midori_rounds_sub_Sub_7_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_23__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_24__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_24__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_7_rs2[4]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[24]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_rs1[4]), .A2(
        Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_24__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[25]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_rs1[4]), .A2(
        Midori_rounds_sub_Sub_7_S1_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_U2 ( .A(r[17]), 
        .B(r[16]), .Z(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_rs2[5]), .B(Midori_rounds_sub_Sub_7_rs1[3]), 
        .ZN(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_7_rs1[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_U4 ( .A(r[17]), 
        .B(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_U2 ( .A(r[12]), 
        .B(Midori_rounds_sub_Sub_7_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_rs2[4]), .B(Midori_rounds_sub_Sub_7_rs2[5]), 
        .Z(Midori_rounds_sub_Sub_7_S1_F_inst_Inst_26__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_1__Compression2_n2), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_1__Compression2_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_7_S1_F_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_7_S1_F_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result1[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[33]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_0__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_0__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[0]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_0__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_U2 ( .A(r[31]), 
        .B(r[30]), .Z(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_7_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_1__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_U2 ( .A(1'b0), .B(
        r[32]), .Z(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_U1 ( .A(1'b0), 
        .B(r[31]), .ZN(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_3__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_3__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_U2 ( .A(r[33]), 
        .B(r[32]), .Z(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_7_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_4__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[5]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_U2 ( .A(1'b0), .B(
        r[34]), .Z(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_U1 ( .A(1'b0), 
        .B(r[33]), .ZN(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_6__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_6__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[6]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_6__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_7__CF_Inst_U4 ( .A(1'b0), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_7__CF_Inst_n9), .Z(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_7__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_7__CF_Inst_n8), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_7__CF_Inst_n7), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_7__CF_Inst_n9) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_7__CF_Inst_n7) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_7__CF_Inst_U1 ( .A(r[34]), 
        .B(r[35]), .Z(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_7__CF_Inst_n8) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_U4 ( .A(r[35]), 
        .B(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_U2 ( .A(r[30]), 
        .B(Midori_rounds_sub_Sub_7_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_U1 ( .A(1'b0), .B(
        1'b0), .Z(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_8__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_9__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_9__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[9]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[1]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_U1 ( .A(r[18]), 
        .B(r[19]), .Z(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_10__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[11]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_U4 ( .A(r[19]), 
        .B(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_U2 ( .A(r[20]), 
        .B(Midori_rounds_sub_Sub_7_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_12__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[1]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_U1 ( .A(r[20]), 
        .B(r[21]), .Z(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_13__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[14]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_U4 ( .A(r[21]), 
        .B(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_U2 ( .A(r[22]), 
        .B(Midori_rounds_sub_Sub_7_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_15__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_15__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[15]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_U2 ( .A(r[23]), 
        .B(r[22]), .Z(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_7_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_n13), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_n12), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_n12) );
  INV_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[1]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_U2 ( .A(r[23]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_n13)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_U1 ( .A(r[18]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_17__CF_Inst_n15)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_18__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_18__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[18]) );
  AOI21_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_18__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_18__CF_Inst_n6) );
  OAI21_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_18__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_U3 ( .A(r[24]), 
        .B(r[25]), .ZN(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[2]), .B1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[1]), .B2(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_19__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[20]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[1]), .C2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_U1 ( .A(r[26]), 
        .B(r[25]), .Z(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_20__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_21__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_21__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[21]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_21__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_21__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_U3 ( .A(r[26]), 
        .B(r[27]), .ZN(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[2]), .B1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[1]), .B2(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_22__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[23]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_U1 ( .A(r[28]), 
        .B(r[27]), .Z(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_23__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_24__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_24__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[24]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_24__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[25]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[3]), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_n9), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_U1 ( .A(r[28]), 
        .B(r[29]), .ZN(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_25__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Out[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_U4 ( .A(r[24]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_n16)
         );
  XOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_U3 ( .A(r[29]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_n17)
         );
  AOI22_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[2]), .B1(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[32]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[32]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[32]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[34]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[34]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[34]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[35]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[35]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[35]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_7_S1_G_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_7_S1_G_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_InAff_out3_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_S2_InAff_out3[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_InAff_out3_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_S2_InAff_out3[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_InAff_out3_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_S2_InAff_out3[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_InAff_out3_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_7_S2_InAff_out3[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_S2_InAff_out2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_rs2[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_S2_InAff_out2[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_rs2[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_S2_InAff_out2[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_rs2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_7_S2_InAff_out2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_3_), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_S2_InAff_out1[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_rs2[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_S2_InAff_out1[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_rs2[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_S2_InAff_out1[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_rs2[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_7_S2_InAff_out1[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_3_), .QN() );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_InputAffine_U3 ( .A(
        Midori_rounds_sub_Sub_7_S2_InAff_out3[1]), .B(Midori_rounds_n979), .Z(
        Midori_rounds_sub_Sub_7_S2_InAff_out3[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_InputAffine_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_InAff_out2[1]), .B(Midori_rounds_n915), .Z(
        Midori_rounds_sub_Sub_7_S2_InAff_out2[3]) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_InputAffine_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_InAff_out1[1]), .B(Midori_rounds_n851), .Z(
        Midori_rounds_sub_Sub_7_S2_InAff_out1[3]) );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_rs2[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_rs2[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_0__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_rs1[0]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_0__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[0]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_0__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_rs2[1]), .C2(Midori_rounds_sub_Sub_7_rs2[2]), 
        .A(Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_0__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_0__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_rs2[1]), .A2(Midori_rounds_sub_Sub_7_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_0__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_7_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_U3 ( .A(r[36]), 
        .B(r[37]), .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_3_), .B2(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[1]), .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_1__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[2]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_7_rs2[1]), .C2(Midori_rounds_sub_Sub_7_rs2[2]), 
        .A(Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_7_rs2[1]), .A2(Midori_rounds_sub_Sub_7_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_rs1[1]), .B(Midori_rounds_sub_Sub_7_rs1[0]), 
        .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_U1 ( .A(r[38]), 
        .B(r[37]), .Z(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_3__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_rs1[0]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_3__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[3]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_3__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_3__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_3__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_3__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_n16), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_7_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_U3 ( .A(r[38]), 
        .B(r[39]), .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_n14)
         );
  OAI21_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[3]), .B2(
        Midori_rounds_sub_Sub_7_rs2[4]), .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_n16) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_7_rs2[5]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_4__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[5]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_rs1[1]), .B(Midori_rounds_sub_Sub_7_rs1[0]), 
        .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_U1 ( .A(r[40]), 
        .B(r[39]), .Z(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_6__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_rs1[0]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_6__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[6]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_6__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_rs2[4]), .C2(Midori_rounds_sub_Sub_7_rs2[5]), 
        .A(Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_6__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_6__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_rs2[4]), .A2(Midori_rounds_sub_Sub_7_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_6__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[7]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_7_rs2[4]), .C2(Midori_rounds_sub_Sub_7_rs2[5]), 
        .A(Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_rs2[4]), .A2(Midori_rounds_sub_Sub_7_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_7_rs1[1]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_U1 ( .A(r[40]), 
        .B(r[41]), .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_7__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_n21), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_n20), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[8]) );
  OAI21_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_U5 ( .B1(
        Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_3_), .B2(
        Midori_rounds_sub_Sub_7_rs2[1]), .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_n19), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_n20) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_7_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_n19) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_n18), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_n17), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_n21) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_rs1[1]), .B(r[41]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_n17) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_rs1[0]), .B(r[36]), .Z(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_8__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_9__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_rs1[2]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_9__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[9]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_9__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_rs2[1]), .C2(Midori_rounds_sub_Sub_7_rs2[2]), 
        .A(Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_9__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_9__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_rs2[1]), .A2(Midori_rounds_sub_Sub_7_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_9__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_U3 ( .A(r[42]), 
        .B(r[43]), .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_3_), .A2(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[2]), .B1(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[1]), .B2(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_10__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[11]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_7_rs2[1]), .C2(Midori_rounds_sub_Sub_7_rs2[2]), 
        .A(Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_7_rs2[1]), .A2(Midori_rounds_sub_Sub_7_rs2[2]), 
        .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_rs1[3]), .B(Midori_rounds_sub_Sub_7_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_U1 ( .A(r[44]), 
        .B(r[43]), .Z(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_12__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_rs1[2]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_12__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[12]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_12__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[3]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_12__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_12__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_12__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_U3 ( .A(r[44]), 
        .B(r[45]), .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[3]), .A2(
        Midori_rounds_sub_Sub_7_rs2[5]), .B1(Midori_rounds_sub_Sub_7_rs2[4]), 
        .B2(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_13__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[14]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[1]), .C2(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[2]), .A(
        Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_rs1[3]), .B(Midori_rounds_sub_Sub_7_rs1[2]), 
        .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_U1 ( .A(r[46]), 
        .B(r[45]), .Z(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_15__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_rs1[2]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_15__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[15]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_15__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_rs2[4]), .C2(Midori_rounds_sub_Sub_7_rs2[5]), 
        .A(Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_3_), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_15__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_15__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_rs2[4]), .A2(Midori_rounds_sub_Sub_7_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_15__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[16]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_7_rs2[4]), .C2(Midori_rounds_sub_Sub_7_rs2[5]), 
        .A(Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_3_), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_rs2[4]), .A2(Midori_rounds_sub_Sub_7_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_n9), .B(
        Midori_rounds_sub_Sub_7_rs1[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_U1 ( .A(r[46]), 
        .B(r[47]), .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_16__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_U4 ( .A(r[42]), 
        .B(Midori_rounds_sub_Sub_7_rs1[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_n16) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_U3 ( .A(r[47]), 
        .B(Midori_rounds_sub_Sub_7_rs1[3]), .Z(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_n17) );
  AOI22_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_3_), .A2(
        Midori_rounds_sub_Sub_7_rs2[2]), .B1(Midori_rounds_sub_Sub_7_rs2[1]), 
        .B2(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_17__CF_Inst_n15) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_18__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_rs1[4]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_18__CF_Inst_n3), .Z(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[18]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_18__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_rs2[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_18__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_U2 ( .A(r[49]), 
        .B(r[48]), .Z(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_rs1[5]), .B(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_19__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[20]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_7_rs2[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_U4 ( .A(r[49]), 
        .B(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_U2 ( .A(r[50]), 
        .B(Midori_rounds_sub_Sub_7_rs2[0]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_rs1[4]), .B(Midori_rounds_sub_Sub_7_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_20__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_21__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_21__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_7_rs1[4]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[21]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_21__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_rs2[4]), .A2(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_U2 ( .A(r[51]), 
        .B(r[50]), .Z(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_rs1[5]), .B(Midori_rounds_sub_Sub_7_rs2[5]), 
        .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_22__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[23]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_U4 ( .A(r[51]), 
        .B(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_U2 ( .A(r[52]), 
        .B(Midori_rounds_sub_Sub_7_S2_InAff_out3_reg[0]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_rs1[4]), .B(Midori_rounds_sub_Sub_7_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_23__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_24__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_24__CF_Inst_n3), .B(
        Midori_rounds_sub_Sub_7_rs1[4]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[24]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_rs2[4]), .A2(
        Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_24__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[25]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_rs2[4]), .A2(
        Midori_rounds_sub_Sub_7_S2_InAff_out2_reg_3_), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_U2 ( .A(r[53]), 
        .B(r[52]), .Z(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_rs1[5]), .B(Midori_rounds_sub_Sub_7_rs2[3]), 
        .ZN(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Out[26]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_7_rs2[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_InAff_out1_reg_3_), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_U4 ( .A(r[53]), 
        .B(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_U2 ( .A(r[48]), 
        .B(Midori_rounds_sub_Sub_7_rs2[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_rs1[4]), .B(Midori_rounds_sub_Sub_7_rs1[5]), 
        .Z(Midori_rounds_sub_Sub_7_S2_F_inst_Inst_26__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[5]), .ZN(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[8]), .ZN(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[0]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[11]), .ZN(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_1__Compression2_n2), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[14]), .ZN(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_1__Compression2_n2) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[17]), .ZN(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[20]), .ZN(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[23]), .ZN(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[26]), .ZN(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[3]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_7_S2_F_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_7_S2_F_inst_InstXOR_2__Compression3_n3) );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_areg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result3[61]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_areg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result1[61]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_areg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[0]), .CK(clk), .Q(
        Midori_rounds_SR_Result2[61]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_0_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[0]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[0]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_1_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[1]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[1]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_2_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[2]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[2]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_3_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[3]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[3]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_4_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[4]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[4]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_5_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[5]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[5]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_6_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[6]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[6]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_7_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[7]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[7]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_8_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[8]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[8]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_9_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[9]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[9]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_10_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[10]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[10]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_11_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[11]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[11]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_12_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[12]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[12]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_13_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[13]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[13]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_14_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[14]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[14]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_15_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[15]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[15]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_16_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[16]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[16]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_17_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[17]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[17]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_18_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[18]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[18]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_19_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[19]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[19]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_20_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[20]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[20]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_21_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[21]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[21]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_22_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[22]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[22]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_23_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[23]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[23]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_24_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[24]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[24]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_25_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[25]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[25]), .QN() );
  DFF_X1 Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg_reg_26_ ( .D(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[26]), .CK(clk), .Q(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[26]), .QN() );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_0__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_0__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[0]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_0__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_0__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[1]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_U2 ( .A(r[67]), 
        .B(r[66]), .Z(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_7_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_1__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[2]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_U2 ( .A(1'b0), .B(
        r[68]), .Z(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_U1 ( .A(1'b0), 
        .B(r[67]), .ZN(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_2__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_3__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_3__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[3]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_3__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_3__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[4]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_U2 ( .A(r[69]), 
        .B(r[68]), .Z(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_7_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_4__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[5]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_U2 ( .A(1'b0), .B(
        r[70]), .Z(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_U1 ( .A(1'b0), 
        .B(r[69]), .ZN(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_5__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_6__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_6__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[6]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_6__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_6__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_7__CF_Inst_U4 ( .A(1'b0), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_7__CF_Inst_n9), .Z(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[7]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_7__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_7__CF_Inst_n8), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_7__CF_Inst_n7), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_7__CF_Inst_n9) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_7__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_7__CF_Inst_n7) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_7__CF_Inst_U1 ( .A(r[70]), 
        .B(r[71]), .Z(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_7__CF_Inst_n8) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[8]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_U4 ( .A(r[71]), 
        .B(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_U2 ( .A(r[66]), 
        .B(Midori_rounds_sub_Sub_7_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_U1 ( .A(1'b0), .B(
        1'b0), .Z(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_8__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_9__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_9__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[9]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_9__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_9__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[10]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[1]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_U1 ( .A(r[54]), 
        .B(r[55]), .Z(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_10__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[11]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_U4 ( .A(r[55]), 
        .B(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_U2 ( .A(r[56]), 
        .B(Midori_rounds_sub_Sub_7_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_11__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_12__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_12__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[12]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_12__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_12__CF_Inst_n3) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_U5 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_n12), .Z(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[13]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_n11), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_n12) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_n10) );
  INV_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[1]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_U1 ( .A(r[56]), 
        .B(r[57]), .Z(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_13__CF_Inst_n11)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[14]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_U5 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_n14) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_U4 ( .A(r[57]), 
        .B(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_n13), .Z(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_U2 ( .A(r[58]), 
        .B(Midori_rounds_sub_Sub_7_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_U1 ( .A(1'b0), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_14__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_15__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_15__CF_Inst_n3), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[15]) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_15__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_15__CF_Inst_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[16]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_n10), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_n9), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_n9) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_U2 ( .A(r[59]), 
        .B(r[58]), .Z(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_n10)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_U1 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_7_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_16__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[17]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_n13), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_n12), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_n12) );
  INV_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[1]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_n11) );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_U2 ( .A(r[59]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_n13)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_U1 ( .A(r[54]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_17__CF_Inst_n15)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_18__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_18__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[18]) );
  AOI21_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_18__CF_Inst_U2 ( .B1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_18__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_18__CF_Inst_n6) );
  OAI21_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_18__CF_Inst_U1 ( .B1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_18__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[19]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_U3 ( .A(r[60]), 
        .B(r[61]), .ZN(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[3]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[2]), .B1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[1]), .B2(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_19__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[20]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[1]), .C2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[2]), .A(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_U1 ( .A(r[62]), 
        .B(r[61]), .Z(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_20__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_21__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_21__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[21]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_21__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[3]), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_21__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_21__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_21__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_21__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_n14), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[22]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_U4 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_n12), .B(1'b0), 
        .ZN(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_U3 ( .A(r[62]), 
        .B(r[63]), .ZN(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_n12)
         );
  AOI22_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[3]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[2]), .B1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[1]), .B2(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_n14) );
  INV_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_22__CF_Inst_n11) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_n15), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_n14), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[23]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_U5 ( .C1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[1]), .C2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[2]), .A(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_n13), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_n14) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_U4 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out3[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_n13) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_U3 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_U2 ( .A(1'b0), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_n11)
         );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_U1 ( .A(r[64]), 
        .B(r[63]), .Z(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_23__CF_Inst_n12)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_24__CF_Inst_U3 ( .A(1'b0), 
        .B(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_24__CF_Inst_n6), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[24]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_24__CF_Inst_U2 ( .C1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[3]), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_24__CF_Inst_n5), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_24__CF_Inst_n6) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_24__CF_Inst_U1 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_24__CF_Inst_n5) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_n12), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_n11), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[25]) );
  OAI211_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_U4 ( .C1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[1]), .C2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[2]), .A(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[3]), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_n10), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_n11) );
  NAND2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_U3 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[1]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[2]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_n10) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_n9), .B(1'b0), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_n12) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_U1 ( .A(r[64]), 
        .B(r[65]), .ZN(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_25__CF_Inst_n9)
         );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_U6 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_n19), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_n18), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Out[26]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_U5 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_n17), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_n16), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_n18) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_U4 ( .A(r[60]), 
        .B(1'b0), .ZN(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_n16)
         );
  XOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_U3 ( .A(r[65]), 
        .B(1'b0), .Z(Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_n17)
         );
  AOI22_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_U2 ( .A1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[3]), .A2(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[2]), .B1(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out2[1]), .B2(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_n15), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_n19) );
  INV_X1 Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_Q12_1_out1[3]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_Inst_26__CF_Inst_n15) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_0__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_0__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[2]), .ZN(
        Midori_rounds_SR_Result1[60]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_0__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[0]), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[1]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_0__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_0__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_0__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[5]), .ZN(
        Midori_rounds_SR_Result2[60]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_0__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[3]), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[4]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_0__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_0__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_0__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[8]), .ZN(
        Midori_rounds_SR_Result3[60]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_0__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[6]), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[7]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_0__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_1__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_1__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[11]), .ZN(
        Midori_rounds_SR_Result1[62]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_1__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[9]), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[10]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_1__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_1__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_1__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[14]), .ZN(
        Midori_rounds_SR_Result2[62]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_1__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[12]), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[13]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_1__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_1__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_1__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[17]), .ZN(
        Midori_rounds_SR_Result3[62]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_1__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[15]), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[16]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_1__Compression3_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_2__Compression1_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_2__Compression1_n3), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[20]), .ZN(
        Midori_rounds_SR_Result1[63]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_2__Compression1_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[18]), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[19]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_2__Compression1_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_2__Compression2_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_2__Compression2_n3), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[23]), .ZN(
        Midori_rounds_SR_Result2[63]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_2__Compression2_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[21]), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[22]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_2__Compression2_n3) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_2__Compression3_U2 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_2__Compression3_n3), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[26]), .ZN(
        Midori_rounds_SR_Result3[63]) );
  XNOR2_X1 Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_2__Compression3_U1 ( .A(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[24]), .B(
        Midori_rounds_sub_Sub_7_S2_G_inst_CF_Reg[25]), .ZN(
        Midori_rounds_sub_Sub_7_S2_G_inst_InstXOR_2__Compression3_n3) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U24 ( .A(Midori_rounds_mul_input1[61]), .B(
        Midori_rounds_mul1_MC1_n24), .ZN(Midori_rounds_SR_Inv_Result1[21]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U23 ( .A(Midori_rounds_mul_input1[60]), .B(
        Midori_rounds_mul1_MC1_n23), .ZN(Midori_rounds_SR_Inv_Result1[20]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U22 ( .A(Midori_rounds_mul_input1[51]), .B(
        Midori_rounds_mul1_MC1_n22), .ZN(Midori_rounds_SR_Inv_Result1[43]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U21 ( .A(Midori_rounds_mul_input1[50]), .B(
        Midori_rounds_mul1_MC1_n21), .ZN(Midori_rounds_SR_Inv_Result1[42]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U20 ( .A(Midori_rounds_mul_input1[49]), .B(
        Midori_rounds_mul1_MC1_n20), .ZN(Midori_rounds_SR_Inv_Result1[41]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U19 ( .A(Midori_rounds_mul_input1[48]), .B(
        Midori_rounds_mul1_MC1_n19), .ZN(Midori_rounds_SR_Inv_Result1[40]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U18 ( .A(Midori_rounds_mul_input1[55]), .B(
        Midori_rounds_mul1_MC1_n22), .ZN(Midori_rounds_SR_Inv_Result1[3]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U17 ( .A(Midori_rounds_mul_input1[63]), .B(
        Midori_rounds_mul_input1[59]), .ZN(Midori_rounds_mul1_MC1_n22) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U16 ( .A(Midori_rounds_mul_input1[54]), .B(
        Midori_rounds_mul1_MC1_n21), .ZN(Midori_rounds_SR_Inv_Result1[2]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U15 ( .A(Midori_rounds_mul_input1[62]), .B(
        Midori_rounds_mul_input1[58]), .ZN(Midori_rounds_mul1_MC1_n21) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U14 ( .A(Midori_rounds_mul_input1[53]), .B(
        Midori_rounds_mul1_MC1_n20), .ZN(Midori_rounds_SR_Inv_Result1[1]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U13 ( .A(Midori_rounds_mul_input1[57]), .B(
        Midori_rounds_mul_input1[61]), .ZN(Midori_rounds_mul1_MC1_n20) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U12 ( .A(Midori_rounds_mul_input1[59]), .B(
        Midori_rounds_mul1_MC1_n18), .ZN(Midori_rounds_SR_Inv_Result1[63]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U11 ( .A(Midori_rounds_mul_input1[58]), .B(
        Midori_rounds_mul1_MC1_n17), .ZN(Midori_rounds_SR_Inv_Result1[62]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U10 ( .A(Midori_rounds_mul_input1[57]), .B(
        Midori_rounds_mul1_MC1_n24), .ZN(Midori_rounds_SR_Inv_Result1[61]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U9 ( .A(Midori_rounds_mul_input1[49]), .B(
        Midori_rounds_mul_input1[53]), .ZN(Midori_rounds_mul1_MC1_n24) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U8 ( .A(Midori_rounds_mul_input1[56]), .B(
        Midori_rounds_mul1_MC1_n23), .ZN(Midori_rounds_SR_Inv_Result1[60]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U7 ( .A(Midori_rounds_mul_input1[52]), .B(
        Midori_rounds_mul_input1[48]), .ZN(Midori_rounds_mul1_MC1_n23) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U6 ( .A(Midori_rounds_mul_input1[63]), .B(
        Midori_rounds_mul1_MC1_n18), .ZN(Midori_rounds_SR_Inv_Result1[23]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U5 ( .A(Midori_rounds_mul_input1[51]), .B(
        Midori_rounds_mul_input1[55]), .ZN(Midori_rounds_mul1_MC1_n18) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U4 ( .A(Midori_rounds_mul_input1[62]), .B(
        Midori_rounds_mul1_MC1_n17), .ZN(Midori_rounds_SR_Inv_Result1[22]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U3 ( .A(Midori_rounds_mul_input1[50]), .B(
        Midori_rounds_mul_input1[54]), .ZN(Midori_rounds_mul1_MC1_n17) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U2 ( .A(Midori_rounds_mul_input1[52]), .B(
        Midori_rounds_mul1_MC1_n19), .ZN(Midori_rounds_SR_Inv_Result1[0]) );
  XNOR2_X1 Midori_rounds_mul1_MC1_U1 ( .A(Midori_rounds_mul_input1[60]), .B(
        Midori_rounds_mul_input1[56]), .ZN(Midori_rounds_mul1_MC1_n19) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U24 ( .A(Midori_rounds_mul_input1[45]), .B(
        Midori_rounds_mul1_MC2_n24), .ZN(Midori_rounds_SR_Inv_Result1[45]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U23 ( .A(Midori_rounds_mul_input1[44]), .B(
        Midori_rounds_mul1_MC2_n23), .ZN(Midori_rounds_SR_Inv_Result1[44]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U22 ( .A(Midori_rounds_mul_input1[35]), .B(
        Midori_rounds_mul1_MC2_n22), .ZN(Midori_rounds_SR_Inv_Result1[19]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U21 ( .A(Midori_rounds_mul_input1[34]), .B(
        Midori_rounds_mul1_MC2_n21), .ZN(Midori_rounds_SR_Inv_Result1[18]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U20 ( .A(Midori_rounds_mul_input1[33]), .B(
        Midori_rounds_mul1_MC2_n20), .ZN(Midori_rounds_SR_Inv_Result1[17]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U19 ( .A(Midori_rounds_mul_input1[32]), .B(
        Midori_rounds_mul1_MC2_n19), .ZN(Midori_rounds_SR_Inv_Result1[16]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U18 ( .A(Midori_rounds_mul_input1[39]), .B(
        Midori_rounds_mul1_MC2_n22), .ZN(Midori_rounds_SR_Inv_Result1[59]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U17 ( .A(Midori_rounds_mul_input1[47]), .B(
        Midori_rounds_mul_input1[43]), .ZN(Midori_rounds_mul1_MC2_n22) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U16 ( .A(Midori_rounds_mul_input1[38]), .B(
        Midori_rounds_mul1_MC2_n21), .ZN(Midori_rounds_SR_Inv_Result1[58]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U15 ( .A(Midori_rounds_mul_input1[46]), .B(
        Midori_rounds_mul_input1[42]), .ZN(Midori_rounds_mul1_MC2_n21) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U14 ( .A(Midori_rounds_mul_input1[37]), .B(
        Midori_rounds_mul1_MC2_n20), .ZN(Midori_rounds_SR_Inv_Result1[57]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U13 ( .A(Midori_rounds_mul_input1[41]), .B(
        Midori_rounds_mul_input1[45]), .ZN(Midori_rounds_mul1_MC2_n20) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U12 ( .A(Midori_rounds_mul_input1[43]), .B(
        Midori_rounds_mul1_MC2_n18), .ZN(Midori_rounds_SR_Inv_Result1[7]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U11 ( .A(Midori_rounds_mul_input1[42]), .B(
        Midori_rounds_mul1_MC2_n17), .ZN(Midori_rounds_SR_Inv_Result1[6]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U10 ( .A(Midori_rounds_mul_input1[41]), .B(
        Midori_rounds_mul1_MC2_n24), .ZN(Midori_rounds_SR_Inv_Result1[5]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U9 ( .A(Midori_rounds_mul_input1[33]), .B(
        Midori_rounds_mul_input1[37]), .ZN(Midori_rounds_mul1_MC2_n24) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U8 ( .A(Midori_rounds_mul_input1[40]), .B(
        Midori_rounds_mul1_MC2_n23), .ZN(Midori_rounds_SR_Inv_Result1[4]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U7 ( .A(Midori_rounds_mul_input1[36]), .B(
        Midori_rounds_mul_input1[32]), .ZN(Midori_rounds_mul1_MC2_n23) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U6 ( .A(Midori_rounds_mul_input1[47]), .B(
        Midori_rounds_mul1_MC2_n18), .ZN(Midori_rounds_SR_Inv_Result1[47]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U5 ( .A(Midori_rounds_mul_input1[35]), .B(
        Midori_rounds_mul_input1[39]), .ZN(Midori_rounds_mul1_MC2_n18) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U4 ( .A(Midori_rounds_mul_input1[46]), .B(
        Midori_rounds_mul1_MC2_n17), .ZN(Midori_rounds_SR_Inv_Result1[46]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U3 ( .A(Midori_rounds_mul_input1[34]), .B(
        Midori_rounds_mul_input1[38]), .ZN(Midori_rounds_mul1_MC2_n17) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U2 ( .A(Midori_rounds_mul_input1[36]), .B(
        Midori_rounds_mul1_MC2_n19), .ZN(Midori_rounds_SR_Inv_Result1[56]) );
  XNOR2_X1 Midori_rounds_mul1_MC2_U1 ( .A(Midori_rounds_mul_input1[44]), .B(
        Midori_rounds_mul_input1[40]), .ZN(Midori_rounds_mul1_MC2_n19) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U24 ( .A(Midori_rounds_mul_input1[29]), .B(
        Midori_rounds_mul1_MC3_n24), .ZN(Midori_rounds_SR_Inv_Result1[49]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U23 ( .A(Midori_rounds_mul_input1[28]), .B(
        Midori_rounds_mul1_MC3_n23), .ZN(Midori_rounds_SR_Inv_Result1[48]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U22 ( .A(Midori_rounds_mul_input1[19]), .B(
        Midori_rounds_mul1_MC3_n22), .ZN(Midori_rounds_SR_Inv_Result1[15]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U21 ( .A(Midori_rounds_mul_input1[18]), .B(
        Midori_rounds_mul1_MC3_n21), .ZN(Midori_rounds_SR_Inv_Result1[14]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U20 ( .A(Midori_rounds_mul_input1[17]), .B(
        Midori_rounds_mul1_MC3_n20), .ZN(Midori_rounds_SR_Inv_Result1[13]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U19 ( .A(Midori_rounds_mul_input1[16]), .B(
        Midori_rounds_mul1_MC3_n19), .ZN(Midori_rounds_SR_Inv_Result1[12]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U18 ( .A(Midori_rounds_mul_input1[23]), .B(
        Midori_rounds_mul1_MC3_n22), .ZN(Midori_rounds_SR_Inv_Result1[39]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U17 ( .A(Midori_rounds_mul_input1[31]), .B(
        Midori_rounds_mul_input1[27]), .ZN(Midori_rounds_mul1_MC3_n22) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U16 ( .A(Midori_rounds_mul_input1[22]), .B(
        Midori_rounds_mul1_MC3_n21), .ZN(Midori_rounds_SR_Inv_Result1[38]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U15 ( .A(Midori_rounds_mul_input1[30]), .B(
        Midori_rounds_mul_input1[26]), .ZN(Midori_rounds_mul1_MC3_n21) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U14 ( .A(Midori_rounds_mul_input1[21]), .B(
        Midori_rounds_mul1_MC3_n20), .ZN(Midori_rounds_SR_Inv_Result1[37]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U13 ( .A(Midori_rounds_mul_input1[25]), .B(
        Midori_rounds_mul_input1[29]), .ZN(Midori_rounds_mul1_MC3_n20) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U12 ( .A(Midori_rounds_mul_input1[27]), .B(
        Midori_rounds_mul1_MC3_n18), .ZN(Midori_rounds_SR_Inv_Result1[27]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U11 ( .A(Midori_rounds_mul_input1[26]), .B(
        Midori_rounds_mul1_MC3_n17), .ZN(Midori_rounds_SR_Inv_Result1[26]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U10 ( .A(Midori_rounds_mul_input1[25]), .B(
        Midori_rounds_mul1_MC3_n24), .ZN(Midori_rounds_SR_Inv_Result1[25]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U9 ( .A(Midori_rounds_mul_input1[17]), .B(
        Midori_rounds_mul_input1[21]), .ZN(Midori_rounds_mul1_MC3_n24) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U8 ( .A(Midori_rounds_mul_input1[24]), .B(
        Midori_rounds_mul1_MC3_n23), .ZN(Midori_rounds_SR_Inv_Result1[24]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U7 ( .A(Midori_rounds_mul_input1[20]), .B(
        Midori_rounds_mul_input1[16]), .ZN(Midori_rounds_mul1_MC3_n23) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U6 ( .A(Midori_rounds_mul_input1[31]), .B(
        Midori_rounds_mul1_MC3_n18), .ZN(Midori_rounds_SR_Inv_Result1[51]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U5 ( .A(Midori_rounds_mul_input1[19]), .B(
        Midori_rounds_mul_input1[23]), .ZN(Midori_rounds_mul1_MC3_n18) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U4 ( .A(Midori_rounds_mul_input1[30]), .B(
        Midori_rounds_mul1_MC3_n17), .ZN(Midori_rounds_SR_Inv_Result1[50]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U3 ( .A(Midori_rounds_mul_input1[18]), .B(
        Midori_rounds_mul_input1[22]), .ZN(Midori_rounds_mul1_MC3_n17) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U2 ( .A(Midori_rounds_mul_input1[20]), .B(
        Midori_rounds_mul1_MC3_n19), .ZN(Midori_rounds_SR_Inv_Result1[36]) );
  XNOR2_X1 Midori_rounds_mul1_MC3_U1 ( .A(Midori_rounds_mul_input1[28]), .B(
        Midori_rounds_mul_input1[24]), .ZN(Midori_rounds_mul1_MC3_n19) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U24 ( .A(Midori_rounds_mul_input1[13]), .B(
        Midori_rounds_mul1_MC4_n24), .ZN(Midori_rounds_SR_Inv_Result1[9]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U23 ( .A(Midori_rounds_mul_input1[12]), .B(
        Midori_rounds_mul1_MC4_n23), .ZN(Midori_rounds_SR_Inv_Result1[8]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U22 ( .A(Midori_rounds_mul_input1[3]), .B(
        Midori_rounds_mul1_MC4_n22), .ZN(Midori_rounds_SR_Inv_Result1[55]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U21 ( .A(Midori_rounds_mul_input1[2]), .B(
        Midori_rounds_mul1_MC4_n21), .ZN(Midori_rounds_SR_Inv_Result1[54]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U20 ( .A(Midori_rounds_mul_input1[1]), .B(
        Midori_rounds_mul1_MC4_n20), .ZN(Midori_rounds_SR_Inv_Result1[53]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U19 ( .A(Midori_rounds_mul_input1[0]), .B(
        Midori_rounds_mul1_MC4_n19), .ZN(Midori_rounds_SR_Inv_Result1[52]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U18 ( .A(Midori_rounds_mul_input1[7]), .B(
        Midori_rounds_mul1_MC4_n22), .ZN(Midori_rounds_SR_Inv_Result1[31]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U17 ( .A(Midori_rounds_mul_input1[15]), .B(
        Midori_rounds_mul_input1[11]), .ZN(Midori_rounds_mul1_MC4_n22) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U16 ( .A(Midori_rounds_mul_input1[6]), .B(
        Midori_rounds_mul1_MC4_n21), .ZN(Midori_rounds_SR_Inv_Result1[30]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U15 ( .A(Midori_rounds_mul_input1[14]), .B(
        Midori_rounds_mul_input1[10]), .ZN(Midori_rounds_mul1_MC4_n21) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U14 ( .A(Midori_rounds_mul_input1[5]), .B(
        Midori_rounds_mul1_MC4_n20), .ZN(Midori_rounds_SR_Inv_Result1[29]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U13 ( .A(Midori_rounds_mul_input1[9]), .B(
        Midori_rounds_mul_input1[13]), .ZN(Midori_rounds_mul1_MC4_n20) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U12 ( .A(Midori_rounds_mul_input1[11]), .B(
        Midori_rounds_mul1_MC4_n18), .ZN(Midori_rounds_SR_Inv_Result1[35]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U11 ( .A(Midori_rounds_mul_input1[10]), .B(
        Midori_rounds_mul1_MC4_n17), .ZN(Midori_rounds_SR_Inv_Result1[34]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U10 ( .A(Midori_rounds_mul_input1[9]), .B(
        Midori_rounds_mul1_MC4_n24), .ZN(Midori_rounds_SR_Inv_Result1[33]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U9 ( .A(Midori_rounds_mul_input1[1]), .B(
        Midori_rounds_mul_input1[5]), .ZN(Midori_rounds_mul1_MC4_n24) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U8 ( .A(Midori_rounds_mul_input1[8]), .B(
        Midori_rounds_mul1_MC4_n23), .ZN(Midori_rounds_SR_Inv_Result1[32]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U7 ( .A(Midori_rounds_mul_input1[4]), .B(
        Midori_rounds_mul_input1[0]), .ZN(Midori_rounds_mul1_MC4_n23) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U6 ( .A(Midori_rounds_mul_input1[15]), .B(
        Midori_rounds_mul1_MC4_n18), .ZN(Midori_rounds_SR_Inv_Result1[11]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U5 ( .A(Midori_rounds_mul_input1[3]), .B(
        Midori_rounds_mul_input1[7]), .ZN(Midori_rounds_mul1_MC4_n18) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U4 ( .A(Midori_rounds_mul_input1[14]), .B(
        Midori_rounds_mul1_MC4_n17), .ZN(Midori_rounds_SR_Inv_Result1[10]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U3 ( .A(Midori_rounds_mul_input1[2]), .B(
        Midori_rounds_mul_input1[6]), .ZN(Midori_rounds_mul1_MC4_n17) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U2 ( .A(Midori_rounds_mul_input1[4]), .B(
        Midori_rounds_mul1_MC4_n19), .ZN(Midori_rounds_SR_Inv_Result1[28]) );
  XNOR2_X1 Midori_rounds_mul1_MC4_U1 ( .A(Midori_rounds_mul_input1[12]), .B(
        Midori_rounds_mul_input1[8]), .ZN(Midori_rounds_mul1_MC4_n19) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U24 ( .A(Midori_rounds_mul_input2[61]), .B(
        Midori_rounds_mul2_MC1_n24), .ZN(Midori_rounds_SR_Inv_Result2[21]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U23 ( .A(Midori_rounds_mul_input2[60]), .B(
        Midori_rounds_mul2_MC1_n23), .ZN(Midori_rounds_SR_Inv_Result2[20]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U22 ( .A(Midori_rounds_mul_input2[51]), .B(
        Midori_rounds_mul2_MC1_n22), .ZN(Midori_rounds_SR_Inv_Result2[43]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U21 ( .A(Midori_rounds_mul_input2[50]), .B(
        Midori_rounds_mul2_MC1_n21), .ZN(Midori_rounds_SR_Inv_Result2[42]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U20 ( .A(Midori_rounds_mul_input2[49]), .B(
        Midori_rounds_mul2_MC1_n20), .ZN(Midori_rounds_SR_Inv_Result2[41]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U19 ( .A(Midori_rounds_mul_input2[48]), .B(
        Midori_rounds_mul2_MC1_n19), .ZN(Midori_rounds_SR_Inv_Result2[40]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U18 ( .A(Midori_rounds_mul_input2[55]), .B(
        Midori_rounds_mul2_MC1_n22), .ZN(Midori_rounds_SR_Inv_Result2[3]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U17 ( .A(Midori_rounds_mul_input2[63]), .B(
        Midori_rounds_mul_input2[59]), .ZN(Midori_rounds_mul2_MC1_n22) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U16 ( .A(Midori_rounds_mul_input2[54]), .B(
        Midori_rounds_mul2_MC1_n21), .ZN(Midori_rounds_SR_Inv_Result2[2]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U15 ( .A(Midori_rounds_mul_input2[62]), .B(
        Midori_rounds_mul_input2[58]), .ZN(Midori_rounds_mul2_MC1_n21) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U14 ( .A(Midori_rounds_mul_input2[53]), .B(
        Midori_rounds_mul2_MC1_n20), .ZN(Midori_rounds_SR_Inv_Result2[1]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U13 ( .A(Midori_rounds_mul_input2[57]), .B(
        Midori_rounds_mul_input2[61]), .ZN(Midori_rounds_mul2_MC1_n20) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U12 ( .A(Midori_rounds_mul_input2[59]), .B(
        Midori_rounds_mul2_MC1_n18), .ZN(Midori_rounds_SR_Inv_Result2[63]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U11 ( .A(Midori_rounds_mul_input2[58]), .B(
        Midori_rounds_mul2_MC1_n17), .ZN(Midori_rounds_SR_Inv_Result2[62]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U10 ( .A(Midori_rounds_mul_input2[57]), .B(
        Midori_rounds_mul2_MC1_n24), .ZN(Midori_rounds_SR_Inv_Result2[61]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U9 ( .A(Midori_rounds_mul_input2[49]), .B(
        Midori_rounds_mul_input2[53]), .ZN(Midori_rounds_mul2_MC1_n24) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U8 ( .A(Midori_rounds_mul_input2[56]), .B(
        Midori_rounds_mul2_MC1_n23), .ZN(Midori_rounds_SR_Inv_Result2[60]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U7 ( .A(Midori_rounds_mul_input2[52]), .B(
        Midori_rounds_mul_input2[48]), .ZN(Midori_rounds_mul2_MC1_n23) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U6 ( .A(Midori_rounds_mul_input2[63]), .B(
        Midori_rounds_mul2_MC1_n18), .ZN(Midori_rounds_SR_Inv_Result2[23]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U5 ( .A(Midori_rounds_mul_input2[51]), .B(
        Midori_rounds_mul_input2[55]), .ZN(Midori_rounds_mul2_MC1_n18) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U4 ( .A(Midori_rounds_mul_input2[62]), .B(
        Midori_rounds_mul2_MC1_n17), .ZN(Midori_rounds_SR_Inv_Result2[22]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U3 ( .A(Midori_rounds_mul_input2[50]), .B(
        Midori_rounds_mul_input2[54]), .ZN(Midori_rounds_mul2_MC1_n17) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U2 ( .A(Midori_rounds_mul_input2[52]), .B(
        Midori_rounds_mul2_MC1_n19), .ZN(Midori_rounds_SR_Inv_Result2[0]) );
  XNOR2_X1 Midori_rounds_mul2_MC1_U1 ( .A(Midori_rounds_mul_input2[60]), .B(
        Midori_rounds_mul_input2[56]), .ZN(Midori_rounds_mul2_MC1_n19) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U24 ( .A(Midori_rounds_mul_input2[45]), .B(
        Midori_rounds_mul2_MC2_n24), .ZN(Midori_rounds_SR_Inv_Result2[45]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U23 ( .A(Midori_rounds_mul_input2[44]), .B(
        Midori_rounds_mul2_MC2_n23), .ZN(Midori_rounds_SR_Inv_Result2[44]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U22 ( .A(Midori_rounds_mul_input2[35]), .B(
        Midori_rounds_mul2_MC2_n22), .ZN(Midori_rounds_SR_Inv_Result2[19]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U21 ( .A(Midori_rounds_mul_input2[34]), .B(
        Midori_rounds_mul2_MC2_n21), .ZN(Midori_rounds_SR_Inv_Result2[18]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U20 ( .A(Midori_rounds_mul_input2[33]), .B(
        Midori_rounds_mul2_MC2_n20), .ZN(Midori_rounds_SR_Inv_Result2[17]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U19 ( .A(Midori_rounds_mul_input2[32]), .B(
        Midori_rounds_mul2_MC2_n19), .ZN(Midori_rounds_SR_Inv_Result2[16]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U18 ( .A(Midori_rounds_mul_input2[39]), .B(
        Midori_rounds_mul2_MC2_n22), .ZN(Midori_rounds_SR_Inv_Result2[59]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U17 ( .A(Midori_rounds_mul_input2[47]), .B(
        Midori_rounds_mul_input2[43]), .ZN(Midori_rounds_mul2_MC2_n22) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U16 ( .A(Midori_rounds_mul_input2[38]), .B(
        Midori_rounds_mul2_MC2_n21), .ZN(Midori_rounds_SR_Inv_Result2[58]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U15 ( .A(Midori_rounds_mul_input2[46]), .B(
        Midori_rounds_mul_input2[42]), .ZN(Midori_rounds_mul2_MC2_n21) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U14 ( .A(Midori_rounds_mul_input2[37]), .B(
        Midori_rounds_mul2_MC2_n20), .ZN(Midori_rounds_SR_Inv_Result2[57]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U13 ( .A(Midori_rounds_mul_input2[41]), .B(
        Midori_rounds_mul_input2[45]), .ZN(Midori_rounds_mul2_MC2_n20) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U12 ( .A(Midori_rounds_mul_input2[43]), .B(
        Midori_rounds_mul2_MC2_n18), .ZN(Midori_rounds_SR_Inv_Result2[7]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U11 ( .A(Midori_rounds_mul_input2[42]), .B(
        Midori_rounds_mul2_MC2_n17), .ZN(Midori_rounds_SR_Inv_Result2[6]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U10 ( .A(Midori_rounds_mul_input2[41]), .B(
        Midori_rounds_mul2_MC2_n24), .ZN(Midori_rounds_SR_Inv_Result2[5]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U9 ( .A(Midori_rounds_mul_input2[33]), .B(
        Midori_rounds_mul_input2[37]), .ZN(Midori_rounds_mul2_MC2_n24) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U8 ( .A(Midori_rounds_mul_input2[40]), .B(
        Midori_rounds_mul2_MC2_n23), .ZN(Midori_rounds_SR_Inv_Result2[4]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U7 ( .A(Midori_rounds_mul_input2[36]), .B(
        Midori_rounds_mul_input2[32]), .ZN(Midori_rounds_mul2_MC2_n23) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U6 ( .A(Midori_rounds_mul_input2[47]), .B(
        Midori_rounds_mul2_MC2_n18), .ZN(Midori_rounds_SR_Inv_Result2[47]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U5 ( .A(Midori_rounds_mul_input2[35]), .B(
        Midori_rounds_mul_input2[39]), .ZN(Midori_rounds_mul2_MC2_n18) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U4 ( .A(Midori_rounds_mul_input2[46]), .B(
        Midori_rounds_mul2_MC2_n17), .ZN(Midori_rounds_SR_Inv_Result2[46]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U3 ( .A(Midori_rounds_mul_input2[34]), .B(
        Midori_rounds_mul_input2[38]), .ZN(Midori_rounds_mul2_MC2_n17) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U2 ( .A(Midori_rounds_mul_input2[36]), .B(
        Midori_rounds_mul2_MC2_n19), .ZN(Midori_rounds_SR_Inv_Result2[56]) );
  XNOR2_X1 Midori_rounds_mul2_MC2_U1 ( .A(Midori_rounds_mul_input2[44]), .B(
        Midori_rounds_mul_input2[40]), .ZN(Midori_rounds_mul2_MC2_n19) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U24 ( .A(Midori_rounds_mul_input2[29]), .B(
        Midori_rounds_mul2_MC3_n24), .ZN(Midori_rounds_SR_Inv_Result2[49]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U23 ( .A(Midori_rounds_mul_input2[28]), .B(
        Midori_rounds_mul2_MC3_n23), .ZN(Midori_rounds_SR_Inv_Result2[48]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U22 ( .A(Midori_rounds_mul_input2[19]), .B(
        Midori_rounds_mul2_MC3_n22), .ZN(Midori_rounds_SR_Inv_Result2[15]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U21 ( .A(Midori_rounds_mul_input2[18]), .B(
        Midori_rounds_mul2_MC3_n21), .ZN(Midori_rounds_SR_Inv_Result2[14]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U20 ( .A(Midori_rounds_mul_input2[17]), .B(
        Midori_rounds_mul2_MC3_n20), .ZN(Midori_rounds_SR_Inv_Result2[13]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U19 ( .A(Midori_rounds_mul_input2[16]), .B(
        Midori_rounds_mul2_MC3_n19), .ZN(Midori_rounds_SR_Inv_Result2[12]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U18 ( .A(Midori_rounds_mul_input2[23]), .B(
        Midori_rounds_mul2_MC3_n22), .ZN(Midori_rounds_SR_Inv_Result2[39]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U17 ( .A(Midori_rounds_mul_input2[31]), .B(
        Midori_rounds_mul_input2[27]), .ZN(Midori_rounds_mul2_MC3_n22) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U16 ( .A(Midori_rounds_mul_input2[22]), .B(
        Midori_rounds_mul2_MC3_n21), .ZN(Midori_rounds_SR_Inv_Result2[38]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U15 ( .A(Midori_rounds_mul_input2[30]), .B(
        Midori_rounds_mul_input2[26]), .ZN(Midori_rounds_mul2_MC3_n21) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U14 ( .A(Midori_rounds_mul_input2[21]), .B(
        Midori_rounds_mul2_MC3_n20), .ZN(Midori_rounds_SR_Inv_Result2[37]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U13 ( .A(Midori_rounds_mul_input2[25]), .B(
        Midori_rounds_mul_input2[29]), .ZN(Midori_rounds_mul2_MC3_n20) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U12 ( .A(Midori_rounds_mul_input2[27]), .B(
        Midori_rounds_mul2_MC3_n18), .ZN(Midori_rounds_SR_Inv_Result2[27]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U11 ( .A(Midori_rounds_mul_input2[26]), .B(
        Midori_rounds_mul2_MC3_n17), .ZN(Midori_rounds_SR_Inv_Result2[26]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U10 ( .A(Midori_rounds_mul_input2[25]), .B(
        Midori_rounds_mul2_MC3_n24), .ZN(Midori_rounds_SR_Inv_Result2[25]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U9 ( .A(Midori_rounds_mul_input2[17]), .B(
        Midori_rounds_mul_input2[21]), .ZN(Midori_rounds_mul2_MC3_n24) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U8 ( .A(Midori_rounds_mul_input2[24]), .B(
        Midori_rounds_mul2_MC3_n23), .ZN(Midori_rounds_SR_Inv_Result2[24]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U7 ( .A(Midori_rounds_mul_input2[20]), .B(
        Midori_rounds_mul_input2[16]), .ZN(Midori_rounds_mul2_MC3_n23) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U6 ( .A(Midori_rounds_mul_input2[31]), .B(
        Midori_rounds_mul2_MC3_n18), .ZN(Midori_rounds_SR_Inv_Result2[51]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U5 ( .A(Midori_rounds_mul_input2[19]), .B(
        Midori_rounds_mul_input2[23]), .ZN(Midori_rounds_mul2_MC3_n18) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U4 ( .A(Midori_rounds_mul_input2[30]), .B(
        Midori_rounds_mul2_MC3_n17), .ZN(Midori_rounds_SR_Inv_Result2[50]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U3 ( .A(Midori_rounds_mul_input2[18]), .B(
        Midori_rounds_mul_input2[22]), .ZN(Midori_rounds_mul2_MC3_n17) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U2 ( .A(Midori_rounds_mul_input2[20]), .B(
        Midori_rounds_mul2_MC3_n19), .ZN(Midori_rounds_SR_Inv_Result2[36]) );
  XNOR2_X1 Midori_rounds_mul2_MC3_U1 ( .A(Midori_rounds_mul_input2[28]), .B(
        Midori_rounds_mul_input2[24]), .ZN(Midori_rounds_mul2_MC3_n19) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U24 ( .A(Midori_rounds_mul_input2[13]), .B(
        Midori_rounds_mul2_MC4_n24), .ZN(Midori_rounds_SR_Inv_Result2[9]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U23 ( .A(Midori_rounds_mul_input2[12]), .B(
        Midori_rounds_mul2_MC4_n23), .ZN(Midori_rounds_SR_Inv_Result2[8]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U22 ( .A(Midori_rounds_mul_input2[3]), .B(
        Midori_rounds_mul2_MC4_n22), .ZN(Midori_rounds_SR_Inv_Result2[55]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U21 ( .A(Midori_rounds_mul_input2[2]), .B(
        Midori_rounds_mul2_MC4_n21), .ZN(Midori_rounds_SR_Inv_Result2[54]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U20 ( .A(Midori_rounds_mul_input2[1]), .B(
        Midori_rounds_mul2_MC4_n20), .ZN(Midori_rounds_SR_Inv_Result2[53]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U19 ( .A(Midori_rounds_mul_input2[0]), .B(
        Midori_rounds_mul2_MC4_n19), .ZN(Midori_rounds_SR_Inv_Result2[52]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U18 ( .A(Midori_rounds_mul_input2[7]), .B(
        Midori_rounds_mul2_MC4_n22), .ZN(Midori_rounds_SR_Inv_Result2[31]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U17 ( .A(Midori_rounds_mul_input2[15]), .B(
        Midori_rounds_mul_input2[11]), .ZN(Midori_rounds_mul2_MC4_n22) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U16 ( .A(Midori_rounds_mul_input2[6]), .B(
        Midori_rounds_mul2_MC4_n21), .ZN(Midori_rounds_SR_Inv_Result2[30]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U15 ( .A(Midori_rounds_mul_input2[14]), .B(
        Midori_rounds_mul_input2[10]), .ZN(Midori_rounds_mul2_MC4_n21) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U14 ( .A(Midori_rounds_mul_input2[5]), .B(
        Midori_rounds_mul2_MC4_n20), .ZN(Midori_rounds_SR_Inv_Result2[29]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U13 ( .A(Midori_rounds_mul_input2[9]), .B(
        Midori_rounds_mul_input2[13]), .ZN(Midori_rounds_mul2_MC4_n20) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U12 ( .A(Midori_rounds_mul_input2[11]), .B(
        Midori_rounds_mul2_MC4_n18), .ZN(Midori_rounds_SR_Inv_Result2[35]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U11 ( .A(Midori_rounds_mul_input2[10]), .B(
        Midori_rounds_mul2_MC4_n17), .ZN(Midori_rounds_SR_Inv_Result2[34]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U10 ( .A(Midori_rounds_mul_input2[9]), .B(
        Midori_rounds_mul2_MC4_n24), .ZN(Midori_rounds_SR_Inv_Result2[33]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U9 ( .A(Midori_rounds_mul_input2[1]), .B(
        Midori_rounds_mul_input2[5]), .ZN(Midori_rounds_mul2_MC4_n24) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U8 ( .A(Midori_rounds_mul_input2[8]), .B(
        Midori_rounds_mul2_MC4_n23), .ZN(Midori_rounds_SR_Inv_Result2[32]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U7 ( .A(Midori_rounds_mul_input2[4]), .B(
        Midori_rounds_mul_input2[0]), .ZN(Midori_rounds_mul2_MC4_n23) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U6 ( .A(Midori_rounds_mul_input2[15]), .B(
        Midori_rounds_mul2_MC4_n18), .ZN(Midori_rounds_SR_Inv_Result2[11]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U5 ( .A(Midori_rounds_mul_input2[3]), .B(
        Midori_rounds_mul_input2[7]), .ZN(Midori_rounds_mul2_MC4_n18) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U4 ( .A(Midori_rounds_mul_input2[14]), .B(
        Midori_rounds_mul2_MC4_n17), .ZN(Midori_rounds_SR_Inv_Result2[10]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U3 ( .A(Midori_rounds_mul_input2[2]), .B(
        Midori_rounds_mul_input2[6]), .ZN(Midori_rounds_mul2_MC4_n17) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U2 ( .A(Midori_rounds_mul_input2[4]), .B(
        Midori_rounds_mul2_MC4_n19), .ZN(Midori_rounds_SR_Inv_Result2[28]) );
  XNOR2_X1 Midori_rounds_mul2_MC4_U1 ( .A(Midori_rounds_mul_input2[12]), .B(
        Midori_rounds_mul_input2[8]), .ZN(Midori_rounds_mul2_MC4_n19) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U24 ( .A(Midori_rounds_mul_input3[61]), .B(
        Midori_rounds_mul3_MC1_n24), .ZN(Midori_rounds_SR_Inv_Result3[21]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U23 ( .A(Midori_rounds_mul_input3[60]), .B(
        Midori_rounds_mul3_MC1_n23), .ZN(Midori_rounds_SR_Inv_Result3[20]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U22 ( .A(Midori_rounds_mul_input3[51]), .B(
        Midori_rounds_mul3_MC1_n22), .ZN(Midori_rounds_SR_Inv_Result3[43]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U21 ( .A(Midori_rounds_mul_input3[50]), .B(
        Midori_rounds_mul3_MC1_n21), .ZN(Midori_rounds_SR_Inv_Result3[42]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U20 ( .A(Midori_rounds_mul_input3[49]), .B(
        Midori_rounds_mul3_MC1_n20), .ZN(Midori_rounds_SR_Inv_Result3[41]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U19 ( .A(Midori_rounds_mul_input3[48]), .B(
        Midori_rounds_mul3_MC1_n19), .ZN(Midori_rounds_SR_Inv_Result3[40]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U18 ( .A(Midori_rounds_mul_input3[55]), .B(
        Midori_rounds_mul3_MC1_n22), .ZN(Midori_rounds_SR_Inv_Result3[3]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U17 ( .A(Midori_rounds_mul_input3[63]), .B(
        Midori_rounds_mul_input3[59]), .ZN(Midori_rounds_mul3_MC1_n22) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U16 ( .A(Midori_rounds_mul_input3[54]), .B(
        Midori_rounds_mul3_MC1_n21), .ZN(Midori_rounds_SR_Inv_Result3[2]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U15 ( .A(Midori_rounds_mul_input3[62]), .B(
        Midori_rounds_mul_input3[58]), .ZN(Midori_rounds_mul3_MC1_n21) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U14 ( .A(Midori_rounds_mul_input3[53]), .B(
        Midori_rounds_mul3_MC1_n20), .ZN(Midori_rounds_SR_Inv_Result3[1]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U13 ( .A(Midori_rounds_mul_input3[57]), .B(
        Midori_rounds_mul_input3[61]), .ZN(Midori_rounds_mul3_MC1_n20) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U12 ( .A(Midori_rounds_mul_input3[59]), .B(
        Midori_rounds_mul3_MC1_n18), .ZN(Midori_rounds_SR_Inv_Result3[63]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U11 ( .A(Midori_rounds_mul_input3[58]), .B(
        Midori_rounds_mul3_MC1_n17), .ZN(Midori_rounds_SR_Inv_Result3[62]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U10 ( .A(Midori_rounds_mul_input3[57]), .B(
        Midori_rounds_mul3_MC1_n24), .ZN(Midori_rounds_SR_Inv_Result3[61]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U9 ( .A(Midori_rounds_mul_input3[49]), .B(
        Midori_rounds_mul_input3[53]), .ZN(Midori_rounds_mul3_MC1_n24) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U8 ( .A(Midori_rounds_mul_input3[56]), .B(
        Midori_rounds_mul3_MC1_n23), .ZN(Midori_rounds_SR_Inv_Result3[60]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U7 ( .A(Midori_rounds_mul_input3[52]), .B(
        Midori_rounds_mul_input3[48]), .ZN(Midori_rounds_mul3_MC1_n23) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U6 ( .A(Midori_rounds_mul_input3[63]), .B(
        Midori_rounds_mul3_MC1_n18), .ZN(Midori_rounds_SR_Inv_Result3[23]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U5 ( .A(Midori_rounds_mul_input3[51]), .B(
        Midori_rounds_mul_input3[55]), .ZN(Midori_rounds_mul3_MC1_n18) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U4 ( .A(Midori_rounds_mul_input3[62]), .B(
        Midori_rounds_mul3_MC1_n17), .ZN(Midori_rounds_SR_Inv_Result3[22]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U3 ( .A(Midori_rounds_mul_input3[50]), .B(
        Midori_rounds_mul_input3[54]), .ZN(Midori_rounds_mul3_MC1_n17) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U2 ( .A(Midori_rounds_mul_input3[52]), .B(
        Midori_rounds_mul3_MC1_n19), .ZN(Midori_rounds_SR_Inv_Result3[0]) );
  XNOR2_X1 Midori_rounds_mul3_MC1_U1 ( .A(Midori_rounds_mul_input3[60]), .B(
        Midori_rounds_mul_input3[56]), .ZN(Midori_rounds_mul3_MC1_n19) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U24 ( .A(Midori_rounds_mul_input3[45]), .B(
        Midori_rounds_mul3_MC2_n24), .ZN(Midori_rounds_SR_Inv_Result3[45]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U23 ( .A(Midori_rounds_mul_input3[44]), .B(
        Midori_rounds_mul3_MC2_n23), .ZN(Midori_rounds_SR_Inv_Result3[44]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U22 ( .A(Midori_rounds_mul_input3[35]), .B(
        Midori_rounds_mul3_MC2_n22), .ZN(Midori_rounds_SR_Inv_Result3[19]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U21 ( .A(Midori_rounds_mul_input3[34]), .B(
        Midori_rounds_mul3_MC2_n21), .ZN(Midori_rounds_SR_Inv_Result3[18]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U20 ( .A(Midori_rounds_mul_input3[33]), .B(
        Midori_rounds_mul3_MC2_n20), .ZN(Midori_rounds_SR_Inv_Result3[17]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U19 ( .A(Midori_rounds_mul_input3[32]), .B(
        Midori_rounds_mul3_MC2_n19), .ZN(Midori_rounds_SR_Inv_Result3[16]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U18 ( .A(Midori_rounds_mul_input3[39]), .B(
        Midori_rounds_mul3_MC2_n22), .ZN(Midori_rounds_SR_Inv_Result3[59]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U17 ( .A(Midori_rounds_mul_input3[47]), .B(
        Midori_rounds_mul_input3[43]), .ZN(Midori_rounds_mul3_MC2_n22) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U16 ( .A(Midori_rounds_mul_input3[38]), .B(
        Midori_rounds_mul3_MC2_n21), .ZN(Midori_rounds_SR_Inv_Result3[58]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U15 ( .A(Midori_rounds_mul_input3[46]), .B(
        Midori_rounds_mul_input3[42]), .ZN(Midori_rounds_mul3_MC2_n21) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U14 ( .A(Midori_rounds_mul_input3[37]), .B(
        Midori_rounds_mul3_MC2_n20), .ZN(Midori_rounds_SR_Inv_Result3[57]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U13 ( .A(Midori_rounds_mul_input3[41]), .B(
        Midori_rounds_mul_input3[45]), .ZN(Midori_rounds_mul3_MC2_n20) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U12 ( .A(Midori_rounds_mul_input3[43]), .B(
        Midori_rounds_mul3_MC2_n18), .ZN(Midori_rounds_SR_Inv_Result3[7]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U11 ( .A(Midori_rounds_mul_input3[42]), .B(
        Midori_rounds_mul3_MC2_n17), .ZN(Midori_rounds_SR_Inv_Result3[6]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U10 ( .A(Midori_rounds_mul_input3[41]), .B(
        Midori_rounds_mul3_MC2_n24), .ZN(Midori_rounds_SR_Inv_Result3[5]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U9 ( .A(Midori_rounds_mul_input3[33]), .B(
        Midori_rounds_mul_input3[37]), .ZN(Midori_rounds_mul3_MC2_n24) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U8 ( .A(Midori_rounds_mul_input3[40]), .B(
        Midori_rounds_mul3_MC2_n23), .ZN(Midori_rounds_SR_Inv_Result3[4]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U7 ( .A(Midori_rounds_mul_input3[36]), .B(
        Midori_rounds_mul_input3[32]), .ZN(Midori_rounds_mul3_MC2_n23) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U6 ( .A(Midori_rounds_mul_input3[47]), .B(
        Midori_rounds_mul3_MC2_n18), .ZN(Midori_rounds_SR_Inv_Result3[47]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U5 ( .A(Midori_rounds_mul_input3[35]), .B(
        Midori_rounds_mul_input3[39]), .ZN(Midori_rounds_mul3_MC2_n18) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U4 ( .A(Midori_rounds_mul_input3[46]), .B(
        Midori_rounds_mul3_MC2_n17), .ZN(Midori_rounds_SR_Inv_Result3[46]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U3 ( .A(Midori_rounds_mul_input3[34]), .B(
        Midori_rounds_mul_input3[38]), .ZN(Midori_rounds_mul3_MC2_n17) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U2 ( .A(Midori_rounds_mul_input3[36]), .B(
        Midori_rounds_mul3_MC2_n19), .ZN(Midori_rounds_SR_Inv_Result3[56]) );
  XNOR2_X1 Midori_rounds_mul3_MC2_U1 ( .A(Midori_rounds_mul_input3[44]), .B(
        Midori_rounds_mul_input3[40]), .ZN(Midori_rounds_mul3_MC2_n19) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U24 ( .A(Midori_rounds_mul_input3[29]), .B(
        Midori_rounds_mul3_MC3_n24), .ZN(Midori_rounds_SR_Inv_Result3[49]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U23 ( .A(Midori_rounds_mul_input3[28]), .B(
        Midori_rounds_mul3_MC3_n23), .ZN(Midori_rounds_SR_Inv_Result3[48]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U22 ( .A(Midori_rounds_mul_input3[19]), .B(
        Midori_rounds_mul3_MC3_n22), .ZN(Midori_rounds_SR_Inv_Result3[15]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U21 ( .A(Midori_rounds_mul_input3[18]), .B(
        Midori_rounds_mul3_MC3_n21), .ZN(Midori_rounds_SR_Inv_Result3[14]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U20 ( .A(Midori_rounds_mul_input3[17]), .B(
        Midori_rounds_mul3_MC3_n20), .ZN(Midori_rounds_SR_Inv_Result3[13]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U19 ( .A(Midori_rounds_mul_input3[16]), .B(
        Midori_rounds_mul3_MC3_n19), .ZN(Midori_rounds_SR_Inv_Result3[12]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U18 ( .A(Midori_rounds_mul_input3[23]), .B(
        Midori_rounds_mul3_MC3_n22), .ZN(Midori_rounds_SR_Inv_Result3[39]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U17 ( .A(Midori_rounds_mul_input3[31]), .B(
        Midori_rounds_mul_input3[27]), .ZN(Midori_rounds_mul3_MC3_n22) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U16 ( .A(Midori_rounds_mul_input3[22]), .B(
        Midori_rounds_mul3_MC3_n21), .ZN(Midori_rounds_SR_Inv_Result3[38]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U15 ( .A(Midori_rounds_mul_input3[30]), .B(
        Midori_rounds_mul_input3[26]), .ZN(Midori_rounds_mul3_MC3_n21) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U14 ( .A(Midori_rounds_mul_input3[21]), .B(
        Midori_rounds_mul3_MC3_n20), .ZN(Midori_rounds_SR_Inv_Result3[37]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U13 ( .A(Midori_rounds_mul_input3[25]), .B(
        Midori_rounds_mul_input3[29]), .ZN(Midori_rounds_mul3_MC3_n20) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U12 ( .A(Midori_rounds_mul_input3[27]), .B(
        Midori_rounds_mul3_MC3_n18), .ZN(Midori_rounds_SR_Inv_Result3[27]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U11 ( .A(Midori_rounds_mul_input3[26]), .B(
        Midori_rounds_mul3_MC3_n17), .ZN(Midori_rounds_SR_Inv_Result3[26]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U10 ( .A(Midori_rounds_mul_input3[25]), .B(
        Midori_rounds_mul3_MC3_n24), .ZN(Midori_rounds_SR_Inv_Result3[25]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U9 ( .A(Midori_rounds_mul_input3[17]), .B(
        Midori_rounds_mul_input3[21]), .ZN(Midori_rounds_mul3_MC3_n24) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U8 ( .A(Midori_rounds_mul_input3[24]), .B(
        Midori_rounds_mul3_MC3_n23), .ZN(Midori_rounds_SR_Inv_Result3[24]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U7 ( .A(Midori_rounds_mul_input3[20]), .B(
        Midori_rounds_mul_input3[16]), .ZN(Midori_rounds_mul3_MC3_n23) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U6 ( .A(Midori_rounds_mul_input3[31]), .B(
        Midori_rounds_mul3_MC3_n18), .ZN(Midori_rounds_SR_Inv_Result3[51]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U5 ( .A(Midori_rounds_mul_input3[19]), .B(
        Midori_rounds_mul_input3[23]), .ZN(Midori_rounds_mul3_MC3_n18) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U4 ( .A(Midori_rounds_mul_input3[30]), .B(
        Midori_rounds_mul3_MC3_n17), .ZN(Midori_rounds_SR_Inv_Result3[50]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U3 ( .A(Midori_rounds_mul_input3[18]), .B(
        Midori_rounds_mul_input3[22]), .ZN(Midori_rounds_mul3_MC3_n17) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U2 ( .A(Midori_rounds_mul_input3[20]), .B(
        Midori_rounds_mul3_MC3_n19), .ZN(Midori_rounds_SR_Inv_Result3[36]) );
  XNOR2_X1 Midori_rounds_mul3_MC3_U1 ( .A(Midori_rounds_mul_input3[28]), .B(
        Midori_rounds_mul_input3[24]), .ZN(Midori_rounds_mul3_MC3_n19) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U24 ( .A(Midori_rounds_mul_input3[13]), .B(
        Midori_rounds_mul3_MC4_n24), .ZN(Midori_rounds_SR_Inv_Result3[9]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U23 ( .A(Midori_rounds_mul_input3[12]), .B(
        Midori_rounds_mul3_MC4_n23), .ZN(Midori_rounds_SR_Inv_Result3[8]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U22 ( .A(Midori_rounds_mul_input3[3]), .B(
        Midori_rounds_mul3_MC4_n22), .ZN(Midori_rounds_SR_Inv_Result3[55]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U21 ( .A(Midori_rounds_mul_input3[2]), .B(
        Midori_rounds_mul3_MC4_n21), .ZN(Midori_rounds_SR_Inv_Result3[54]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U20 ( .A(Midori_rounds_mul_input3[1]), .B(
        Midori_rounds_mul3_MC4_n20), .ZN(Midori_rounds_SR_Inv_Result3[53]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U19 ( .A(Midori_rounds_mul_input3[0]), .B(
        Midori_rounds_mul3_MC4_n19), .ZN(Midori_rounds_SR_Inv_Result3[52]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U18 ( .A(Midori_rounds_mul_input3[7]), .B(
        Midori_rounds_mul3_MC4_n22), .ZN(Midori_rounds_SR_Inv_Result3[31]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U17 ( .A(Midori_rounds_mul_input3[15]), .B(
        Midori_rounds_mul_input3[11]), .ZN(Midori_rounds_mul3_MC4_n22) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U16 ( .A(Midori_rounds_mul_input3[6]), .B(
        Midori_rounds_mul3_MC4_n21), .ZN(Midori_rounds_SR_Inv_Result3[30]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U15 ( .A(Midori_rounds_mul_input3[14]), .B(
        Midori_rounds_mul_input3[10]), .ZN(Midori_rounds_mul3_MC4_n21) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U14 ( .A(Midori_rounds_mul_input3[5]), .B(
        Midori_rounds_mul3_MC4_n20), .ZN(Midori_rounds_SR_Inv_Result3[29]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U13 ( .A(Midori_rounds_mul_input3[9]), .B(
        Midori_rounds_mul_input3[13]), .ZN(Midori_rounds_mul3_MC4_n20) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U12 ( .A(Midori_rounds_mul_input3[11]), .B(
        Midori_rounds_mul3_MC4_n18), .ZN(Midori_rounds_SR_Inv_Result3[35]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U11 ( .A(Midori_rounds_mul_input3[10]), .B(
        Midori_rounds_mul3_MC4_n17), .ZN(Midori_rounds_SR_Inv_Result3[34]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U10 ( .A(Midori_rounds_mul_input3[9]), .B(
        Midori_rounds_mul3_MC4_n24), .ZN(Midori_rounds_SR_Inv_Result3[33]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U9 ( .A(Midori_rounds_mul_input3[1]), .B(
        Midori_rounds_mul_input3[5]), .ZN(Midori_rounds_mul3_MC4_n24) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U8 ( .A(Midori_rounds_mul_input3[8]), .B(
        Midori_rounds_mul3_MC4_n23), .ZN(Midori_rounds_SR_Inv_Result3[32]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U7 ( .A(Midori_rounds_mul_input3[4]), .B(
        Midori_rounds_mul_input3[0]), .ZN(Midori_rounds_mul3_MC4_n23) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U6 ( .A(Midori_rounds_mul_input3[15]), .B(
        Midori_rounds_mul3_MC4_n18), .ZN(Midori_rounds_SR_Inv_Result3[11]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U5 ( .A(Midori_rounds_mul_input3[3]), .B(
        Midori_rounds_mul_input3[7]), .ZN(Midori_rounds_mul3_MC4_n18) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U4 ( .A(Midori_rounds_mul_input3[14]), .B(
        Midori_rounds_mul3_MC4_n17), .ZN(Midori_rounds_SR_Inv_Result3[10]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U3 ( .A(Midori_rounds_mul_input3[2]), .B(
        Midori_rounds_mul_input3[6]), .ZN(Midori_rounds_mul3_MC4_n17) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U2 ( .A(Midori_rounds_mul_input3[4]), .B(
        Midori_rounds_mul3_MC4_n19), .ZN(Midori_rounds_SR_Inv_Result3[28]) );
  XNOR2_X1 Midori_rounds_mul3_MC4_U1 ( .A(Midori_rounds_mul_input3[12]), .B(
        Midori_rounds_mul_input3[8]), .ZN(Midori_rounds_mul3_MC4_n19) );
endmodule

