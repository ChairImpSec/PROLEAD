module circuit ( X_s0, X_s1, X_s1_bar, Fresh, reset, clk, Y_s0, Y_s1 );
  input [7:0] X_s0;
  input [7:0] X_s1;
  input [7:0] X_s1_bar;
  input [33:0] Fresh;
  output [7:0] Y_s0;
  output [7:0] Y_s1;
  input reset, clk;
  wire   top_L29, top_new_AGEMA_signal_409, top_new_AGEMA_signal_410, top_L28,
         top_new_AGEMA_signal_407, top_new_AGEMA_signal_408, top_L27,
         top_new_AGEMA_signal_405, top_new_AGEMA_signal_406, top_L26,
         top_new_AGEMA_signal_403, top_new_AGEMA_signal_404, top_L25,
         top_new_AGEMA_signal_401, top_new_AGEMA_signal_402, top_L24,
         top_new_AGEMA_signal_399, top_new_AGEMA_signal_400, top_L23,
         top_new_AGEMA_signal_389, top_new_AGEMA_signal_390, top_L22,
         top_new_AGEMA_signal_387, top_new_AGEMA_signal_388, top_L21,
         top_new_AGEMA_signal_397, top_new_AGEMA_signal_398, top_L20,
         top_new_AGEMA_signal_395, top_new_AGEMA_signal_396, top_L19,
         top_new_AGEMA_signal_385, top_new_AGEMA_signal_386, top_L18,
         top_new_AGEMA_signal_371, top_new_AGEMA_signal_372, top_L17,
         top_new_AGEMA_signal_369, top_new_AGEMA_signal_370, top_L16,
         top_new_AGEMA_signal_393, top_new_AGEMA_signal_394, top_L15,
         top_new_AGEMA_signal_367, top_new_AGEMA_signal_368, top_L14,
         top_new_AGEMA_signal_365, top_new_AGEMA_signal_366, top_L13,
         top_new_AGEMA_signal_391, top_new_AGEMA_signal_392, top_L12,
         top_new_AGEMA_signal_351, top_new_AGEMA_signal_352, top_L11,
         top_new_AGEMA_signal_383, top_new_AGEMA_signal_384, top_L10,
         top_new_AGEMA_signal_381, top_new_AGEMA_signal_382, top_L9,
         top_new_AGEMA_signal_379, top_new_AGEMA_signal_380, top_L8,
         top_new_AGEMA_signal_349, top_new_AGEMA_signal_350, top_L7,
         top_new_AGEMA_signal_377, top_new_AGEMA_signal_378, top_L6,
         top_new_AGEMA_signal_375, top_new_AGEMA_signal_376, top_L5,
         top_new_AGEMA_signal_363, top_new_AGEMA_signal_364, top_L4,
         top_new_AGEMA_signal_361, top_new_AGEMA_signal_362, top_L3,
         top_new_AGEMA_signal_359, top_new_AGEMA_signal_360, top_L2,
         top_new_AGEMA_signal_357, top_new_AGEMA_signal_358, top_L1,
         top_new_AGEMA_signal_347, top_new_AGEMA_signal_348, top_L0,
         top_new_AGEMA_signal_373, top_new_AGEMA_signal_374,
         top_new_AGEMA_signal_345, top_new_AGEMA_signal_346,
         top_new_AGEMA_signal_355, top_new_AGEMA_signal_356,
         top_new_AGEMA_signal_343, top_new_AGEMA_signal_344,
         top_new_AGEMA_signal_327, top_new_AGEMA_signal_328,
         top_new_AGEMA_signal_325, top_new_AGEMA_signal_326,
         top_new_AGEMA_signal_341, top_new_AGEMA_signal_342,
         top_new_AGEMA_signal_323, top_new_AGEMA_signal_324,
         top_new_AGEMA_signal_321, top_new_AGEMA_signal_322,
         top_new_AGEMA_signal_339, top_new_AGEMA_signal_340,
         top_new_AGEMA_signal_337, top_new_AGEMA_signal_338,
         top_new_AGEMA_signal_353, top_new_AGEMA_signal_354,
         top_new_AGEMA_signal_335, top_new_AGEMA_signal_336,
         top_new_AGEMA_signal_319, top_new_AGEMA_signal_320,
         top_new_AGEMA_signal_317, top_new_AGEMA_signal_318,
         top_new_AGEMA_signal_333, top_new_AGEMA_signal_334,
         top_new_AGEMA_signal_315, top_new_AGEMA_signal_316,
         top_new_AGEMA_signal_313, top_new_AGEMA_signal_314,
         top_new_AGEMA_signal_331, top_new_AGEMA_signal_332, top_M45,
         top_new_AGEMA_signal_329, top_new_AGEMA_signal_330, top_M44,
         top_new_AGEMA_signal_311, top_new_AGEMA_signal_312, top_M43,
         top_new_AGEMA_signal_309, top_new_AGEMA_signal_310, top_M42,
         top_new_AGEMA_signal_307, top_new_AGEMA_signal_308, top_M41,
         top_new_AGEMA_signal_305, top_new_AGEMA_signal_306, top_M40,
         top_new_AGEMA_signal_303, top_new_AGEMA_signal_304, top_M39,
         top_new_AGEMA_signal_301, top_new_AGEMA_signal_302, top_M38,
         top_new_AGEMA_signal_299, top_new_AGEMA_signal_300, top_M37,
         top_new_AGEMA_signal_297, top_new_AGEMA_signal_298, top_M36,
         top_new_AGEMA_signal_295, top_new_AGEMA_signal_296,
         top_new_AGEMA_signal_293, top_new_AGEMA_signal_294,
         top_new_AGEMA_signal_275, top_new_AGEMA_signal_276, top_M33,
         top_new_AGEMA_signal_285, top_new_AGEMA_signal_286,
         top_new_AGEMA_signal_291, top_new_AGEMA_signal_292,
         top_new_AGEMA_signal_283, top_new_AGEMA_signal_284,
         top_new_AGEMA_signal_289, top_new_AGEMA_signal_290,
         top_new_AGEMA_signal_287, top_new_AGEMA_signal_288, top_M28,
         top_new_AGEMA_signal_281, top_new_AGEMA_signal_282, top_M27,
         top_new_AGEMA_signal_273, top_new_AGEMA_signal_274, top_M26,
         top_new_AGEMA_signal_279, top_new_AGEMA_signal_280,
         top_new_AGEMA_signal_271, top_new_AGEMA_signal_272, top_M24,
         top_new_AGEMA_signal_277, top_new_AGEMA_signal_278, top_M23,
         top_new_AGEMA_signal_269, top_new_AGEMA_signal_270, top_M22,
         top_new_AGEMA_signal_267, top_new_AGEMA_signal_268, top_M21,
         top_new_AGEMA_signal_265, top_new_AGEMA_signal_266, top_M20,
         top_new_AGEMA_signal_263, top_new_AGEMA_signal_264, top_M19,
         top_new_AGEMA_signal_261, top_new_AGEMA_signal_262, top_M18,
         top_new_AGEMA_signal_259, top_new_AGEMA_signal_260, top_M17,
         top_new_AGEMA_signal_257, top_new_AGEMA_signal_258, top_M16,
         top_new_AGEMA_signal_255, top_new_AGEMA_signal_256, top_M15,
         top_new_AGEMA_signal_253, top_new_AGEMA_signal_254,
         top_new_AGEMA_signal_249, top_new_AGEMA_signal_250, top_M13,
         top_new_AGEMA_signal_247, top_new_AGEMA_signal_248,
         top_new_AGEMA_signal_231, top_new_AGEMA_signal_232,
         top_new_AGEMA_signal_229, top_new_AGEMA_signal_230, top_M10,
         top_new_AGEMA_signal_251, top_new_AGEMA_signal_252,
         top_new_AGEMA_signal_245, top_new_AGEMA_signal_246, top_M8,
         top_new_AGEMA_signal_243, top_new_AGEMA_signal_244,
         top_new_AGEMA_signal_227, top_new_AGEMA_signal_228,
         top_new_AGEMA_signal_225, top_new_AGEMA_signal_226, top_M5,
         top_new_AGEMA_signal_241, top_new_AGEMA_signal_242,
         top_new_AGEMA_signal_223, top_new_AGEMA_signal_224, top_M3,
         top_new_AGEMA_signal_239, top_new_AGEMA_signal_240,
         top_new_AGEMA_signal_237, top_new_AGEMA_signal_238,
         top_new_AGEMA_signal_221, top_new_AGEMA_signal_222, top_T27,
         top_new_AGEMA_signal_205, top_new_AGEMA_signal_206, top_T26,
         top_new_AGEMA_signal_219, top_new_AGEMA_signal_220, top_T25,
         top_new_AGEMA_signal_235, top_new_AGEMA_signal_236, top_T24,
         top_new_AGEMA_signal_233, top_new_AGEMA_signal_234, top_T23,
         top_new_AGEMA_signal_217, top_new_AGEMA_signal_218, top_T22,
         top_new_AGEMA_signal_203, top_new_AGEMA_signal_204, top_T21,
         top_new_AGEMA_signal_189, top_new_AGEMA_signal_190, top_T20,
         top_new_AGEMA_signal_215, top_new_AGEMA_signal_216, top_T19,
         top_new_AGEMA_signal_201, top_new_AGEMA_signal_202, top_T18,
         top_new_AGEMA_signal_187, top_new_AGEMA_signal_188, top_T17,
         top_new_AGEMA_signal_213, top_new_AGEMA_signal_214, top_T16,
         top_new_AGEMA_signal_199, top_new_AGEMA_signal_200, top_T15,
         top_new_AGEMA_signal_197, top_new_AGEMA_signal_198, top_T14,
         top_new_AGEMA_signal_211, top_new_AGEMA_signal_212, top_T13,
         top_new_AGEMA_signal_195, top_new_AGEMA_signal_196, top_T12,
         top_new_AGEMA_signal_183, top_new_AGEMA_signal_184, top_T11,
         top_new_AGEMA_signal_181, top_new_AGEMA_signal_182, top_T10,
         top_new_AGEMA_signal_209, top_new_AGEMA_signal_210, top_T9,
         top_new_AGEMA_signal_193, top_new_AGEMA_signal_194, top_T8,
         top_new_AGEMA_signal_207, top_new_AGEMA_signal_208, top_T7,
         top_new_AGEMA_signal_179, top_new_AGEMA_signal_180, top_T6,
         top_new_AGEMA_signal_191, top_new_AGEMA_signal_192, top_T5,
         top_new_AGEMA_signal_173, top_new_AGEMA_signal_174, top_T4,
         top_new_AGEMA_signal_169, top_new_AGEMA_signal_170, top_T3,
         top_new_AGEMA_signal_167, top_new_AGEMA_signal_168, top_T2,
         top_new_AGEMA_signal_163, top_new_AGEMA_signal_164, top_T1,
         top_new_AGEMA_signal_159, top_new_AGEMA_signal_160,
         top_XOR_T1_U1_xorInst_n4, top_XOR_T1_U1_xorInst_n3,
         top_XOR_T1_U1_xorInst_n2, top_XOR_T1_U1_xorInst_n1,
         top_XOR_T2_U1_xorInst_n12, top_XOR_T2_U1_xorInst_n11,
         top_XOR_T2_U1_xorInst_n10, top_XOR_T2_U1_xorInst_n9,
         top_XOR_T3_U1_xorInst_n12, top_XOR_T3_U1_xorInst_n11,
         top_XOR_T3_U1_xorInst_n10, top_XOR_T3_U1_xorInst_n9,
         top_XOR_T4_U1_xorInst_n12, top_XOR_T4_U1_xorInst_n11,
         top_XOR_T4_U1_xorInst_n10, top_XOR_T4_U1_xorInst_n9,
         top_XOR_T5_U1_xorInst_n12, top_XOR_T5_U1_xorInst_n11,
         top_XOR_T5_U1_xorInst_n10, top_XOR_T5_U1_xorInst_n9,
         top_XOR_T6_U1_xorInst_n12, top_XOR_T6_U1_xorInst_n11,
         top_XOR_T6_U1_xorInst_n10, top_XOR_T6_U1_xorInst_n9,
         top_XOR_T7_U1_xorInst_n12, top_XOR_T7_U1_xorInst_n11,
         top_XOR_T7_U1_xorInst_n10, top_XOR_T7_U1_xorInst_n9,
         top_XOR_T8_U1_xorInst_n12, top_XOR_T8_U1_xorInst_n11,
         top_XOR_T8_U1_xorInst_n10, top_XOR_T8_U1_xorInst_n9,
         top_XOR_T9_U1_xorInst_n12, top_XOR_T9_U1_xorInst_n11,
         top_XOR_T9_U1_xorInst_n10, top_XOR_T9_U1_xorInst_n9,
         top_XOR_T10_U1_xorInst_n12, top_XOR_T10_U1_xorInst_n11,
         top_XOR_T10_U1_xorInst_n10, top_XOR_T10_U1_xorInst_n9,
         top_XOR_T11_U1_xorInst_n12, top_XOR_T11_U1_xorInst_n11,
         top_XOR_T11_U1_xorInst_n10, top_XOR_T11_U1_xorInst_n9,
         top_XOR_T12_U1_xorInst_n12, top_XOR_T12_U1_xorInst_n11,
         top_XOR_T12_U1_xorInst_n10, top_XOR_T12_U1_xorInst_n9,
         top_XOR_T13_U1_xorInst_n12, top_XOR_T13_U1_xorInst_n11,
         top_XOR_T13_U1_xorInst_n10, top_XOR_T13_U1_xorInst_n9,
         top_XOR_T14_U1_xorInst_n12, top_XOR_T14_U1_xorInst_n11,
         top_XOR_T14_U1_xorInst_n10, top_XOR_T14_U1_xorInst_n9,
         top_XOR_T15_U1_xorInst_n12, top_XOR_T15_U1_xorInst_n11,
         top_XOR_T15_U1_xorInst_n10, top_XOR_T15_U1_xorInst_n9,
         top_XOR_T16_U1_xorInst_n12, top_XOR_T16_U1_xorInst_n11,
         top_XOR_T16_U1_xorInst_n10, top_XOR_T16_U1_xorInst_n9,
         top_XOR_T17_U1_xorInst_n12, top_XOR_T17_U1_xorInst_n11,
         top_XOR_T17_U1_xorInst_n10, top_XOR_T17_U1_xorInst_n9,
         top_XOR_T18_U1_xorInst_n12, top_XOR_T18_U1_xorInst_n11,
         top_XOR_T18_U1_xorInst_n10, top_XOR_T18_U1_xorInst_n9,
         top_XOR_T19_U1_xorInst_n12, top_XOR_T19_U1_xorInst_n11,
         top_XOR_T19_U1_xorInst_n10, top_XOR_T19_U1_xorInst_n9,
         top_XOR_T20_U1_xorInst_n12, top_XOR_T20_U1_xorInst_n11,
         top_XOR_T20_U1_xorInst_n10, top_XOR_T20_U1_xorInst_n9,
         top_XOR_T21_U1_xorInst_n12, top_XOR_T21_U1_xorInst_n11,
         top_XOR_T21_U1_xorInst_n10, top_XOR_T21_U1_xorInst_n9,
         top_XOR_T22_U1_xorInst_n12, top_XOR_T22_U1_xorInst_n11,
         top_XOR_T22_U1_xorInst_n10, top_XOR_T22_U1_xorInst_n9,
         top_XOR_T23_U1_xorInst_n12, top_XOR_T23_U1_xorInst_n11,
         top_XOR_T23_U1_xorInst_n10, top_XOR_T23_U1_xorInst_n9,
         top_XOR_T24_U1_xorInst_n12, top_XOR_T24_U1_xorInst_n11,
         top_XOR_T24_U1_xorInst_n10, top_XOR_T24_U1_xorInst_n9,
         top_XOR_T25_U1_xorInst_n12, top_XOR_T25_U1_xorInst_n11,
         top_XOR_T25_U1_xorInst_n10, top_XOR_T25_U1_xorInst_n9,
         top_XOR_T26_U1_xorInst_n12, top_XOR_T26_U1_xorInst_n11,
         top_XOR_T26_U1_xorInst_n10, top_XOR_T26_U1_xorInst_n9,
         top_XOR_T27_U1_xorInst_n12, top_XOR_T27_U1_xorInst_n11,
         top_XOR_T27_U1_xorInst_n10, top_XOR_T27_U1_xorInst_n9,
         top_AND_M1_U1_nonlinearInst_n18, top_AND_M1_U1_nonlinearInst_n17,
         top_AND_M1_U1_nonlinearInst_n16, top_AND_M1_U1_nonlinearInst_n15,
         top_AND_M1_U1_nonlinearInst_n14, top_AND_M1_U1_nonlinearInst_n13,
         top_AND_M1_U1_nonlinearInst_n12, top_AND_M1_U1_nonlinearInst_n11,
         top_AND_M1_U1_nonlinearInst_n10, top_AND_M1_U1_nonlinearInst_n9,
         top_AND_M1_U1_nonlinearInst_n8, top_AND_M1_U1_nonlinearInst_n7,
         top_AND_M1_U1_nonlinearInst_n6, top_AND_M1_U1_nonlinearInst_n5,
         top_AND_M1_U1_nonlinearInst_n4, top_AND_M1_U1_nonlinearInst_n3,
         top_AND_M1_U1_nonlinearInst_n2, top_AND_M1_U1_nonlinearInst_n1,
         top_AND_M1_U1_gen_reg_0__regIns_n2,
         top_AND_M1_U1_gen_reg_0__regIns_N3,
         top_AND_M1_U1_gen_reg_1__regIns_n2,
         top_AND_M1_U1_gen_reg_1__regIns_N3,
         top_AND_M1_U1_gen_reg_2__regIns_n2,
         top_AND_M1_U1_gen_reg_2__regIns_N3,
         top_AND_M1_U1_gen_reg_3__regIns_n2,
         top_AND_M1_U1_gen_reg_3__regIns_N3,
         top_AND_M1_U1_gen_reg_4__regIns_n2,
         top_AND_M1_U1_gen_reg_4__regIns_N3,
         top_AND_M1_U1_gen_reg_5__regIns_n2,
         top_AND_M1_U1_gen_reg_5__regIns_N3,
         top_AND_M1_U1_gen_reg_6__regIns_n2,
         top_AND_M1_U1_gen_reg_6__regIns_N3,
         top_AND_M1_U1_gen_reg_7__regIns_n2,
         top_AND_M1_U1_gen_reg_7__regIns_N3,
         top_AND_M1_U1_OperationInst_andInst0_n1,
         top_AND_M1_U1_OperationInst_andInst1_n3,
         top_AND_M1_U1_OperationInst_andInst2_n3,
         top_AND_M1_U1_OperationInst_andInst3_n3,
         top_AND_M1_U1_OperationInst_orInst1_n2,
         top_AND_M1_U1_OperationInst_orInst1_n1,
         top_AND_M1_U1_OperationInst_andInst4_n3,
         top_AND_M1_U1_OperationInst_andInst5_n3,
         top_AND_M1_U1_OperationInst_andInst6_n3,
         top_AND_M1_U1_OperationInst_andInst7_n3,
         top_AND_M1_U1_OperationInst_orInst2_n6,
         top_AND_M1_U1_OperationInst_orInst2_n5,
         top_AND_M2_U1_nonlinearInst_n64, top_AND_M2_U1_nonlinearInst_n63,
         top_AND_M2_U1_nonlinearInst_n62, top_AND_M2_U1_nonlinearInst_n61,
         top_AND_M2_U1_nonlinearInst_n60, top_AND_M2_U1_nonlinearInst_n59,
         top_AND_M2_U1_nonlinearInst_n58, top_AND_M2_U1_nonlinearInst_n57,
         top_AND_M2_U1_nonlinearInst_n56, top_AND_M2_U1_nonlinearInst_n55,
         top_AND_M2_U1_nonlinearInst_n54, top_AND_M2_U1_nonlinearInst_n53,
         top_AND_M2_U1_nonlinearInst_n52, top_AND_M2_U1_nonlinearInst_n51,
         top_AND_M2_U1_nonlinearInst_n50, top_AND_M2_U1_nonlinearInst_n49,
         top_AND_M2_U1_nonlinearInst_n48, top_AND_M2_U1_nonlinearInst_n47,
         top_AND_M2_U1_gen_reg_0__regIns_n2,
         top_AND_M2_U1_gen_reg_0__regIns_N3,
         top_AND_M2_U1_gen_reg_1__regIns_n2,
         top_AND_M2_U1_gen_reg_1__regIns_N3,
         top_AND_M2_U1_gen_reg_2__regIns_n2,
         top_AND_M2_U1_gen_reg_2__regIns_N3,
         top_AND_M2_U1_gen_reg_3__regIns_n2,
         top_AND_M2_U1_gen_reg_3__regIns_N3,
         top_AND_M2_U1_gen_reg_4__regIns_n2,
         top_AND_M2_U1_gen_reg_4__regIns_N3,
         top_AND_M2_U1_gen_reg_5__regIns_n2,
         top_AND_M2_U1_gen_reg_5__regIns_N3,
         top_AND_M2_U1_gen_reg_6__regIns_n2,
         top_AND_M2_U1_gen_reg_6__regIns_N3,
         top_AND_M2_U1_gen_reg_7__regIns_n2,
         top_AND_M2_U1_gen_reg_7__regIns_N3,
         top_AND_M2_U1_OperationInst_andInst0_n3,
         top_AND_M2_U1_OperationInst_andInst1_n3,
         top_AND_M2_U1_OperationInst_andInst2_n3,
         top_AND_M2_U1_OperationInst_andInst3_n3,
         top_AND_M2_U1_OperationInst_orInst1_n6,
         top_AND_M2_U1_OperationInst_orInst1_n5,
         top_AND_M2_U1_OperationInst_andInst4_n3,
         top_AND_M2_U1_OperationInst_andInst5_n3,
         top_AND_M2_U1_OperationInst_andInst6_n3,
         top_AND_M2_U1_OperationInst_andInst7_n3,
         top_AND_M2_U1_OperationInst_orInst2_n6,
         top_AND_M2_U1_OperationInst_orInst2_n5, top_XOR_M3_U1_xorInst_n12,
         top_XOR_M3_U1_xorInst_n11, top_XOR_M3_U1_xorInst_n10,
         top_XOR_M3_U1_xorInst_n9, top_AND_M4_U1_nonlinearInst_n64,
         top_AND_M4_U1_nonlinearInst_n63, top_AND_M4_U1_nonlinearInst_n62,
         top_AND_M4_U1_nonlinearInst_n61, top_AND_M4_U1_nonlinearInst_n60,
         top_AND_M4_U1_nonlinearInst_n59, top_AND_M4_U1_nonlinearInst_n58,
         top_AND_M4_U1_nonlinearInst_n57, top_AND_M4_U1_nonlinearInst_n56,
         top_AND_M4_U1_nonlinearInst_n55, top_AND_M4_U1_nonlinearInst_n54,
         top_AND_M4_U1_nonlinearInst_n53, top_AND_M4_U1_nonlinearInst_n52,
         top_AND_M4_U1_nonlinearInst_n51, top_AND_M4_U1_nonlinearInst_n50,
         top_AND_M4_U1_nonlinearInst_n49, top_AND_M4_U1_nonlinearInst_n48,
         top_AND_M4_U1_nonlinearInst_n47, top_AND_M4_U1_gen_reg_0__regIns_n2,
         top_AND_M4_U1_gen_reg_0__regIns_N3,
         top_AND_M4_U1_gen_reg_1__regIns_n2,
         top_AND_M4_U1_gen_reg_1__regIns_N3,
         top_AND_M4_U1_gen_reg_2__regIns_n2,
         top_AND_M4_U1_gen_reg_2__regIns_N3,
         top_AND_M4_U1_gen_reg_3__regIns_n2,
         top_AND_M4_U1_gen_reg_3__regIns_N3,
         top_AND_M4_U1_gen_reg_4__regIns_n2,
         top_AND_M4_U1_gen_reg_4__regIns_N3,
         top_AND_M4_U1_gen_reg_5__regIns_n2,
         top_AND_M4_U1_gen_reg_5__regIns_N3,
         top_AND_M4_U1_gen_reg_6__regIns_n2,
         top_AND_M4_U1_gen_reg_6__regIns_N3,
         top_AND_M4_U1_gen_reg_7__regIns_n2,
         top_AND_M4_U1_gen_reg_7__regIns_N3,
         top_AND_M4_U1_OperationInst_andInst0_n3,
         top_AND_M4_U1_OperationInst_andInst1_n3,
         top_AND_M4_U1_OperationInst_andInst2_n3,
         top_AND_M4_U1_OperationInst_andInst3_n3,
         top_AND_M4_U1_OperationInst_orInst1_n6,
         top_AND_M4_U1_OperationInst_orInst1_n5,
         top_AND_M4_U1_OperationInst_andInst4_n3,
         top_AND_M4_U1_OperationInst_andInst5_n3,
         top_AND_M4_U1_OperationInst_andInst6_n3,
         top_AND_M4_U1_OperationInst_andInst7_n3,
         top_AND_M4_U1_OperationInst_orInst2_n6,
         top_AND_M4_U1_OperationInst_orInst2_n5, top_XOR_M5_U1_xorInst_n12,
         top_XOR_M5_U1_xorInst_n11, top_XOR_M5_U1_xorInst_n10,
         top_XOR_M5_U1_xorInst_n9, top_AND_M6_U1_nonlinearInst_n64,
         top_AND_M6_U1_nonlinearInst_n63, top_AND_M6_U1_nonlinearInst_n62,
         top_AND_M6_U1_nonlinearInst_n61, top_AND_M6_U1_nonlinearInst_n60,
         top_AND_M6_U1_nonlinearInst_n59, top_AND_M6_U1_nonlinearInst_n58,
         top_AND_M6_U1_nonlinearInst_n57, top_AND_M6_U1_nonlinearInst_n56,
         top_AND_M6_U1_nonlinearInst_n55, top_AND_M6_U1_nonlinearInst_n54,
         top_AND_M6_U1_nonlinearInst_n53, top_AND_M6_U1_nonlinearInst_n52,
         top_AND_M6_U1_nonlinearInst_n51, top_AND_M6_U1_nonlinearInst_n50,
         top_AND_M6_U1_nonlinearInst_n49, top_AND_M6_U1_nonlinearInst_n48,
         top_AND_M6_U1_nonlinearInst_n47, top_AND_M6_U1_gen_reg_0__regIns_n2,
         top_AND_M6_U1_gen_reg_0__regIns_N3,
         top_AND_M6_U1_gen_reg_1__regIns_n2,
         top_AND_M6_U1_gen_reg_1__regIns_N3,
         top_AND_M6_U1_gen_reg_2__regIns_n2,
         top_AND_M6_U1_gen_reg_2__regIns_N3,
         top_AND_M6_U1_gen_reg_3__regIns_n2,
         top_AND_M6_U1_gen_reg_3__regIns_N3,
         top_AND_M6_U1_gen_reg_4__regIns_n2,
         top_AND_M6_U1_gen_reg_4__regIns_N3,
         top_AND_M6_U1_gen_reg_5__regIns_n2,
         top_AND_M6_U1_gen_reg_5__regIns_N3,
         top_AND_M6_U1_gen_reg_6__regIns_n2,
         top_AND_M6_U1_gen_reg_6__regIns_N3,
         top_AND_M6_U1_gen_reg_7__regIns_n2,
         top_AND_M6_U1_gen_reg_7__regIns_N3,
         top_AND_M6_U1_OperationInst_andInst0_n3,
         top_AND_M6_U1_OperationInst_andInst1_n3,
         top_AND_M6_U1_OperationInst_andInst2_n3,
         top_AND_M6_U1_OperationInst_andInst3_n3,
         top_AND_M6_U1_OperationInst_orInst1_n6,
         top_AND_M6_U1_OperationInst_orInst1_n5,
         top_AND_M6_U1_OperationInst_andInst4_n3,
         top_AND_M6_U1_OperationInst_andInst5_n3,
         top_AND_M6_U1_OperationInst_andInst6_n3,
         top_AND_M6_U1_OperationInst_andInst7_n3,
         top_AND_M6_U1_OperationInst_orInst2_n6,
         top_AND_M6_U1_OperationInst_orInst2_n5,
         top_AND_M7_U1_nonlinearInst_n64, top_AND_M7_U1_nonlinearInst_n63,
         top_AND_M7_U1_nonlinearInst_n62, top_AND_M7_U1_nonlinearInst_n61,
         top_AND_M7_U1_nonlinearInst_n60, top_AND_M7_U1_nonlinearInst_n59,
         top_AND_M7_U1_nonlinearInst_n58, top_AND_M7_U1_nonlinearInst_n57,
         top_AND_M7_U1_nonlinearInst_n56, top_AND_M7_U1_nonlinearInst_n55,
         top_AND_M7_U1_nonlinearInst_n54, top_AND_M7_U1_nonlinearInst_n53,
         top_AND_M7_U1_nonlinearInst_n52, top_AND_M7_U1_nonlinearInst_n51,
         top_AND_M7_U1_nonlinearInst_n50, top_AND_M7_U1_nonlinearInst_n49,
         top_AND_M7_U1_nonlinearInst_n48, top_AND_M7_U1_nonlinearInst_n47,
         top_AND_M7_U1_gen_reg_0__regIns_n2,
         top_AND_M7_U1_gen_reg_0__regIns_N3,
         top_AND_M7_U1_gen_reg_1__regIns_n2,
         top_AND_M7_U1_gen_reg_1__regIns_N3,
         top_AND_M7_U1_gen_reg_2__regIns_n2,
         top_AND_M7_U1_gen_reg_2__regIns_N3,
         top_AND_M7_U1_gen_reg_3__regIns_n2,
         top_AND_M7_U1_gen_reg_3__regIns_N3,
         top_AND_M7_U1_gen_reg_4__regIns_n2,
         top_AND_M7_U1_gen_reg_4__regIns_N3,
         top_AND_M7_U1_gen_reg_5__regIns_n2,
         top_AND_M7_U1_gen_reg_5__regIns_N3,
         top_AND_M7_U1_gen_reg_6__regIns_n2,
         top_AND_M7_U1_gen_reg_6__regIns_N3,
         top_AND_M7_U1_gen_reg_7__regIns_n2,
         top_AND_M7_U1_gen_reg_7__regIns_N3,
         top_AND_M7_U1_OperationInst_andInst0_n3,
         top_AND_M7_U1_OperationInst_andInst1_n3,
         top_AND_M7_U1_OperationInst_andInst2_n3,
         top_AND_M7_U1_OperationInst_andInst3_n3,
         top_AND_M7_U1_OperationInst_orInst1_n6,
         top_AND_M7_U1_OperationInst_orInst1_n5,
         top_AND_M7_U1_OperationInst_andInst4_n3,
         top_AND_M7_U1_OperationInst_andInst5_n3,
         top_AND_M7_U1_OperationInst_andInst6_n3,
         top_AND_M7_U1_OperationInst_andInst7_n3,
         top_AND_M7_U1_OperationInst_orInst2_n6,
         top_AND_M7_U1_OperationInst_orInst2_n5, top_XOR_M8_U1_xorInst_n12,
         top_XOR_M8_U1_xorInst_n11, top_XOR_M8_U1_xorInst_n10,
         top_XOR_M8_U1_xorInst_n9, top_AND_M9_U1_nonlinearInst_n64,
         top_AND_M9_U1_nonlinearInst_n63, top_AND_M9_U1_nonlinearInst_n62,
         top_AND_M9_U1_nonlinearInst_n61, top_AND_M9_U1_nonlinearInst_n60,
         top_AND_M9_U1_nonlinearInst_n59, top_AND_M9_U1_nonlinearInst_n58,
         top_AND_M9_U1_nonlinearInst_n57, top_AND_M9_U1_nonlinearInst_n56,
         top_AND_M9_U1_nonlinearInst_n55, top_AND_M9_U1_nonlinearInst_n54,
         top_AND_M9_U1_nonlinearInst_n53, top_AND_M9_U1_nonlinearInst_n52,
         top_AND_M9_U1_nonlinearInst_n51, top_AND_M9_U1_nonlinearInst_n50,
         top_AND_M9_U1_nonlinearInst_n49, top_AND_M9_U1_nonlinearInst_n48,
         top_AND_M9_U1_nonlinearInst_n47, top_AND_M9_U1_gen_reg_0__regIns_n2,
         top_AND_M9_U1_gen_reg_0__regIns_N3,
         top_AND_M9_U1_gen_reg_1__regIns_n2,
         top_AND_M9_U1_gen_reg_1__regIns_N3,
         top_AND_M9_U1_gen_reg_2__regIns_n2,
         top_AND_M9_U1_gen_reg_2__regIns_N3,
         top_AND_M9_U1_gen_reg_3__regIns_n2,
         top_AND_M9_U1_gen_reg_3__regIns_N3,
         top_AND_M9_U1_gen_reg_4__regIns_n2,
         top_AND_M9_U1_gen_reg_4__regIns_N3,
         top_AND_M9_U1_gen_reg_5__regIns_n2,
         top_AND_M9_U1_gen_reg_5__regIns_N3,
         top_AND_M9_U1_gen_reg_6__regIns_n2,
         top_AND_M9_U1_gen_reg_6__regIns_N3,
         top_AND_M9_U1_gen_reg_7__regIns_n2,
         top_AND_M9_U1_gen_reg_7__regIns_N3,
         top_AND_M9_U1_OperationInst_andInst0_n3,
         top_AND_M9_U1_OperationInst_andInst1_n3,
         top_AND_M9_U1_OperationInst_andInst2_n3,
         top_AND_M9_U1_OperationInst_andInst3_n3,
         top_AND_M9_U1_OperationInst_orInst1_n6,
         top_AND_M9_U1_OperationInst_orInst1_n5,
         top_AND_M9_U1_OperationInst_andInst4_n3,
         top_AND_M9_U1_OperationInst_andInst5_n3,
         top_AND_M9_U1_OperationInst_andInst6_n3,
         top_AND_M9_U1_OperationInst_andInst7_n3,
         top_AND_M9_U1_OperationInst_orInst2_n6,
         top_AND_M9_U1_OperationInst_orInst2_n5, top_XOR_M10_U1_xorInst_n12,
         top_XOR_M10_U1_xorInst_n11, top_XOR_M10_U1_xorInst_n10,
         top_XOR_M10_U1_xorInst_n9, top_AND_M11_U1_nonlinearInst_n64,
         top_AND_M11_U1_nonlinearInst_n63, top_AND_M11_U1_nonlinearInst_n62,
         top_AND_M11_U1_nonlinearInst_n61, top_AND_M11_U1_nonlinearInst_n60,
         top_AND_M11_U1_nonlinearInst_n59, top_AND_M11_U1_nonlinearInst_n58,
         top_AND_M11_U1_nonlinearInst_n57, top_AND_M11_U1_nonlinearInst_n56,
         top_AND_M11_U1_nonlinearInst_n55, top_AND_M11_U1_nonlinearInst_n54,
         top_AND_M11_U1_nonlinearInst_n53, top_AND_M11_U1_nonlinearInst_n52,
         top_AND_M11_U1_nonlinearInst_n51, top_AND_M11_U1_nonlinearInst_n50,
         top_AND_M11_U1_nonlinearInst_n49, top_AND_M11_U1_nonlinearInst_n48,
         top_AND_M11_U1_nonlinearInst_n47, top_AND_M11_U1_gen_reg_0__regIns_n2,
         top_AND_M11_U1_gen_reg_0__regIns_N3,
         top_AND_M11_U1_gen_reg_1__regIns_n2,
         top_AND_M11_U1_gen_reg_1__regIns_N3,
         top_AND_M11_U1_gen_reg_2__regIns_n2,
         top_AND_M11_U1_gen_reg_2__regIns_N3,
         top_AND_M11_U1_gen_reg_3__regIns_n2,
         top_AND_M11_U1_gen_reg_3__regIns_N3,
         top_AND_M11_U1_gen_reg_4__regIns_n2,
         top_AND_M11_U1_gen_reg_4__regIns_N3,
         top_AND_M11_U1_gen_reg_5__regIns_n2,
         top_AND_M11_U1_gen_reg_5__regIns_N3,
         top_AND_M11_U1_gen_reg_6__regIns_n2,
         top_AND_M11_U1_gen_reg_6__regIns_N3,
         top_AND_M11_U1_gen_reg_7__regIns_n2,
         top_AND_M11_U1_gen_reg_7__regIns_N3,
         top_AND_M11_U1_OperationInst_andInst0_n3,
         top_AND_M11_U1_OperationInst_andInst1_n3,
         top_AND_M11_U1_OperationInst_andInst2_n3,
         top_AND_M11_U1_OperationInst_andInst3_n3,
         top_AND_M11_U1_OperationInst_orInst1_n6,
         top_AND_M11_U1_OperationInst_orInst1_n5,
         top_AND_M11_U1_OperationInst_andInst4_n3,
         top_AND_M11_U1_OperationInst_andInst5_n3,
         top_AND_M11_U1_OperationInst_andInst6_n3,
         top_AND_M11_U1_OperationInst_andInst7_n3,
         top_AND_M11_U1_OperationInst_orInst2_n6,
         top_AND_M11_U1_OperationInst_orInst2_n5,
         top_AND_M12_U1_nonlinearInst_n64, top_AND_M12_U1_nonlinearInst_n63,
         top_AND_M12_U1_nonlinearInst_n62, top_AND_M12_U1_nonlinearInst_n61,
         top_AND_M12_U1_nonlinearInst_n60, top_AND_M12_U1_nonlinearInst_n59,
         top_AND_M12_U1_nonlinearInst_n58, top_AND_M12_U1_nonlinearInst_n57,
         top_AND_M12_U1_nonlinearInst_n56, top_AND_M12_U1_nonlinearInst_n55,
         top_AND_M12_U1_nonlinearInst_n54, top_AND_M12_U1_nonlinearInst_n53,
         top_AND_M12_U1_nonlinearInst_n52, top_AND_M12_U1_nonlinearInst_n51,
         top_AND_M12_U1_nonlinearInst_n50, top_AND_M12_U1_nonlinearInst_n49,
         top_AND_M12_U1_nonlinearInst_n48, top_AND_M12_U1_nonlinearInst_n47,
         top_AND_M12_U1_gen_reg_0__regIns_n2,
         top_AND_M12_U1_gen_reg_0__regIns_N3,
         top_AND_M12_U1_gen_reg_1__regIns_n2,
         top_AND_M12_U1_gen_reg_1__regIns_N3,
         top_AND_M12_U1_gen_reg_2__regIns_n2,
         top_AND_M12_U1_gen_reg_2__regIns_N3,
         top_AND_M12_U1_gen_reg_3__regIns_n2,
         top_AND_M12_U1_gen_reg_3__regIns_N3,
         top_AND_M12_U1_gen_reg_4__regIns_n2,
         top_AND_M12_U1_gen_reg_4__regIns_N3,
         top_AND_M12_U1_gen_reg_5__regIns_n2,
         top_AND_M12_U1_gen_reg_5__regIns_N3,
         top_AND_M12_U1_gen_reg_6__regIns_n2,
         top_AND_M12_U1_gen_reg_6__regIns_N3,
         top_AND_M12_U1_gen_reg_7__regIns_n2,
         top_AND_M12_U1_gen_reg_7__regIns_N3,
         top_AND_M12_U1_OperationInst_andInst0_n3,
         top_AND_M12_U1_OperationInst_andInst1_n3,
         top_AND_M12_U1_OperationInst_andInst2_n3,
         top_AND_M12_U1_OperationInst_andInst3_n3,
         top_AND_M12_U1_OperationInst_orInst1_n6,
         top_AND_M12_U1_OperationInst_orInst1_n5,
         top_AND_M12_U1_OperationInst_andInst4_n3,
         top_AND_M12_U1_OperationInst_andInst5_n3,
         top_AND_M12_U1_OperationInst_andInst6_n3,
         top_AND_M12_U1_OperationInst_andInst7_n3,
         top_AND_M12_U1_OperationInst_orInst2_n6,
         top_AND_M12_U1_OperationInst_orInst2_n5, top_XOR_M13_U1_xorInst_n12,
         top_XOR_M13_U1_xorInst_n11, top_XOR_M13_U1_xorInst_n10,
         top_XOR_M13_U1_xorInst_n9, top_AND_M14_U1_nonlinearInst_n64,
         top_AND_M14_U1_nonlinearInst_n63, top_AND_M14_U1_nonlinearInst_n62,
         top_AND_M14_U1_nonlinearInst_n61, top_AND_M14_U1_nonlinearInst_n60,
         top_AND_M14_U1_nonlinearInst_n59, top_AND_M14_U1_nonlinearInst_n58,
         top_AND_M14_U1_nonlinearInst_n57, top_AND_M14_U1_nonlinearInst_n56,
         top_AND_M14_U1_nonlinearInst_n55, top_AND_M14_U1_nonlinearInst_n54,
         top_AND_M14_U1_nonlinearInst_n53, top_AND_M14_U1_nonlinearInst_n52,
         top_AND_M14_U1_nonlinearInst_n51, top_AND_M14_U1_nonlinearInst_n50,
         top_AND_M14_U1_nonlinearInst_n49, top_AND_M14_U1_nonlinearInst_n48,
         top_AND_M14_U1_nonlinearInst_n47, top_AND_M14_U1_gen_reg_0__regIns_n2,
         top_AND_M14_U1_gen_reg_0__regIns_N3,
         top_AND_M14_U1_gen_reg_1__regIns_n2,
         top_AND_M14_U1_gen_reg_1__regIns_N3,
         top_AND_M14_U1_gen_reg_2__regIns_n2,
         top_AND_M14_U1_gen_reg_2__regIns_N3,
         top_AND_M14_U1_gen_reg_3__regIns_n2,
         top_AND_M14_U1_gen_reg_3__regIns_N3,
         top_AND_M14_U1_gen_reg_4__regIns_n2,
         top_AND_M14_U1_gen_reg_4__regIns_N3,
         top_AND_M14_U1_gen_reg_5__regIns_n2,
         top_AND_M14_U1_gen_reg_5__regIns_N3,
         top_AND_M14_U1_gen_reg_6__regIns_n2,
         top_AND_M14_U1_gen_reg_6__regIns_N3,
         top_AND_M14_U1_gen_reg_7__regIns_n2,
         top_AND_M14_U1_gen_reg_7__regIns_N3,
         top_AND_M14_U1_OperationInst_andInst0_n3,
         top_AND_M14_U1_OperationInst_andInst1_n3,
         top_AND_M14_U1_OperationInst_andInst2_n3,
         top_AND_M14_U1_OperationInst_andInst3_n3,
         top_AND_M14_U1_OperationInst_orInst1_n6,
         top_AND_M14_U1_OperationInst_orInst1_n5,
         top_AND_M14_U1_OperationInst_andInst4_n3,
         top_AND_M14_U1_OperationInst_andInst5_n3,
         top_AND_M14_U1_OperationInst_andInst6_n3,
         top_AND_M14_U1_OperationInst_andInst7_n3,
         top_AND_M14_U1_OperationInst_orInst2_n6,
         top_AND_M14_U1_OperationInst_orInst2_n5, top_XOR_M15_U1_xorInst_n12,
         top_XOR_M15_U1_xorInst_n11, top_XOR_M15_U1_xorInst_n10,
         top_XOR_M15_U1_xorInst_n9, top_XOR_M16_U1_xorInst_n12,
         top_XOR_M16_U1_xorInst_n11, top_XOR_M16_U1_xorInst_n10,
         top_XOR_M16_U1_xorInst_n9, top_XOR_M17_U1_xorInst_n12,
         top_XOR_M17_U1_xorInst_n11, top_XOR_M17_U1_xorInst_n10,
         top_XOR_M17_U1_xorInst_n9, top_XOR_M18_U1_xorInst_n12,
         top_XOR_M18_U1_xorInst_n11, top_XOR_M18_U1_xorInst_n10,
         top_XOR_M18_U1_xorInst_n9, top_XOR_M19_U1_xorInst_n12,
         top_XOR_M19_U1_xorInst_n11, top_XOR_M19_U1_xorInst_n10,
         top_XOR_M19_U1_xorInst_n9, top_XOR_M20_U1_xorInst_n12,
         top_XOR_M20_U1_xorInst_n11, top_XOR_M20_U1_xorInst_n10,
         top_XOR_M20_U1_xorInst_n9, top_XOR_M21_U1_xorInst_n12,
         top_XOR_M21_U1_xorInst_n11, top_XOR_M21_U1_xorInst_n10,
         top_XOR_M21_U1_xorInst_n9, top_XOR_M22_U1_xorInst_n12,
         top_XOR_M22_U1_xorInst_n11, top_XOR_M22_U1_xorInst_n10,
         top_XOR_M22_U1_xorInst_n9, top_XOR_M23_U1_xorInst_n12,
         top_XOR_M23_U1_xorInst_n11, top_XOR_M23_U1_xorInst_n10,
         top_XOR_M23_U1_xorInst_n9, top_XOR_M24_U1_xorInst_n12,
         top_XOR_M24_U1_xorInst_n11, top_XOR_M24_U1_xorInst_n10,
         top_XOR_M24_U1_xorInst_n9, top_AND_M25_U1_nonlinearInst_n64,
         top_AND_M25_U1_nonlinearInst_n63, top_AND_M25_U1_nonlinearInst_n62,
         top_AND_M25_U1_nonlinearInst_n61, top_AND_M25_U1_nonlinearInst_n60,
         top_AND_M25_U1_nonlinearInst_n59, top_AND_M25_U1_nonlinearInst_n58,
         top_AND_M25_U1_nonlinearInst_n57, top_AND_M25_U1_nonlinearInst_n56,
         top_AND_M25_U1_nonlinearInst_n55, top_AND_M25_U1_nonlinearInst_n54,
         top_AND_M25_U1_nonlinearInst_n53, top_AND_M25_U1_nonlinearInst_n52,
         top_AND_M25_U1_nonlinearInst_n51, top_AND_M25_U1_nonlinearInst_n50,
         top_AND_M25_U1_nonlinearInst_n49, top_AND_M25_U1_nonlinearInst_n48,
         top_AND_M25_U1_nonlinearInst_n47, top_AND_M25_U1_gen_reg_0__regIns_n2,
         top_AND_M25_U1_gen_reg_0__regIns_N3,
         top_AND_M25_U1_gen_reg_1__regIns_n2,
         top_AND_M25_U1_gen_reg_1__regIns_N3,
         top_AND_M25_U1_gen_reg_2__regIns_n2,
         top_AND_M25_U1_gen_reg_2__regIns_N3,
         top_AND_M25_U1_gen_reg_3__regIns_n2,
         top_AND_M25_U1_gen_reg_3__regIns_N3,
         top_AND_M25_U1_gen_reg_4__regIns_n2,
         top_AND_M25_U1_gen_reg_4__regIns_N3,
         top_AND_M25_U1_gen_reg_5__regIns_n2,
         top_AND_M25_U1_gen_reg_5__regIns_N3,
         top_AND_M25_U1_gen_reg_6__regIns_n2,
         top_AND_M25_U1_gen_reg_6__regIns_N3,
         top_AND_M25_U1_gen_reg_7__regIns_n2,
         top_AND_M25_U1_gen_reg_7__regIns_N3,
         top_AND_M25_U1_OperationInst_andInst0_n3,
         top_AND_M25_U1_OperationInst_andInst1_n3,
         top_AND_M25_U1_OperationInst_andInst2_n3,
         top_AND_M25_U1_OperationInst_andInst3_n3,
         top_AND_M25_U1_OperationInst_orInst1_n6,
         top_AND_M25_U1_OperationInst_orInst1_n5,
         top_AND_M25_U1_OperationInst_andInst4_n3,
         top_AND_M25_U1_OperationInst_andInst5_n3,
         top_AND_M25_U1_OperationInst_andInst6_n3,
         top_AND_M25_U1_OperationInst_andInst7_n3,
         top_AND_M25_U1_OperationInst_orInst2_n6,
         top_AND_M25_U1_OperationInst_orInst2_n5, top_XOR_M26_U1_xorInst_n12,
         top_XOR_M26_U1_xorInst_n11, top_XOR_M26_U1_xorInst_n10,
         top_XOR_M26_U1_xorInst_n9, top_XOR_M27_U1_xorInst_n12,
         top_XOR_M27_U1_xorInst_n11, top_XOR_M27_U1_xorInst_n10,
         top_XOR_M27_U1_xorInst_n9, top_XOR_M28_U1_xorInst_n12,
         top_XOR_M28_U1_xorInst_n11, top_XOR_M28_U1_xorInst_n10,
         top_XOR_M28_U1_xorInst_n9, top_AND_M29_U1_nonlinearInst_n64,
         top_AND_M29_U1_nonlinearInst_n63, top_AND_M29_U1_nonlinearInst_n62,
         top_AND_M29_U1_nonlinearInst_n61, top_AND_M29_U1_nonlinearInst_n60,
         top_AND_M29_U1_nonlinearInst_n59, top_AND_M29_U1_nonlinearInst_n58,
         top_AND_M29_U1_nonlinearInst_n57, top_AND_M29_U1_nonlinearInst_n56,
         top_AND_M29_U1_nonlinearInst_n55, top_AND_M29_U1_nonlinearInst_n54,
         top_AND_M29_U1_nonlinearInst_n53, top_AND_M29_U1_nonlinearInst_n52,
         top_AND_M29_U1_nonlinearInst_n51, top_AND_M29_U1_nonlinearInst_n50,
         top_AND_M29_U1_nonlinearInst_n49, top_AND_M29_U1_nonlinearInst_n48,
         top_AND_M29_U1_nonlinearInst_n47, top_AND_M29_U1_gen_reg_0__regIns_n2,
         top_AND_M29_U1_gen_reg_0__regIns_N3,
         top_AND_M29_U1_gen_reg_1__regIns_n2,
         top_AND_M29_U1_gen_reg_1__regIns_N3,
         top_AND_M29_U1_gen_reg_2__regIns_n2,
         top_AND_M29_U1_gen_reg_2__regIns_N3,
         top_AND_M29_U1_gen_reg_3__regIns_n2,
         top_AND_M29_U1_gen_reg_3__regIns_N3,
         top_AND_M29_U1_gen_reg_4__regIns_n2,
         top_AND_M29_U1_gen_reg_4__regIns_N3,
         top_AND_M29_U1_gen_reg_5__regIns_n2,
         top_AND_M29_U1_gen_reg_5__regIns_N3,
         top_AND_M29_U1_gen_reg_6__regIns_n2,
         top_AND_M29_U1_gen_reg_6__regIns_N3,
         top_AND_M29_U1_gen_reg_7__regIns_n2,
         top_AND_M29_U1_gen_reg_7__regIns_N3,
         top_AND_M29_U1_OperationInst_andInst0_n3,
         top_AND_M29_U1_OperationInst_andInst1_n3,
         top_AND_M29_U1_OperationInst_andInst2_n3,
         top_AND_M29_U1_OperationInst_andInst3_n3,
         top_AND_M29_U1_OperationInst_orInst1_n6,
         top_AND_M29_U1_OperationInst_orInst1_n5,
         top_AND_M29_U1_OperationInst_andInst4_n3,
         top_AND_M29_U1_OperationInst_andInst5_n3,
         top_AND_M29_U1_OperationInst_andInst6_n3,
         top_AND_M29_U1_OperationInst_andInst7_n3,
         top_AND_M29_U1_OperationInst_orInst2_n6,
         top_AND_M29_U1_OperationInst_orInst2_n5,
         top_AND_M30_U1_nonlinearInst_n64, top_AND_M30_U1_nonlinearInst_n63,
         top_AND_M30_U1_nonlinearInst_n62, top_AND_M30_U1_nonlinearInst_n61,
         top_AND_M30_U1_nonlinearInst_n60, top_AND_M30_U1_nonlinearInst_n59,
         top_AND_M30_U1_nonlinearInst_n58, top_AND_M30_U1_nonlinearInst_n57,
         top_AND_M30_U1_nonlinearInst_n56, top_AND_M30_U1_nonlinearInst_n55,
         top_AND_M30_U1_nonlinearInst_n54, top_AND_M30_U1_nonlinearInst_n53,
         top_AND_M30_U1_nonlinearInst_n52, top_AND_M30_U1_nonlinearInst_n51,
         top_AND_M30_U1_nonlinearInst_n50, top_AND_M30_U1_nonlinearInst_n49,
         top_AND_M30_U1_nonlinearInst_n48, top_AND_M30_U1_nonlinearInst_n47,
         top_AND_M30_U1_gen_reg_0__regIns_n2,
         top_AND_M30_U1_gen_reg_0__regIns_N3,
         top_AND_M30_U1_gen_reg_1__regIns_n2,
         top_AND_M30_U1_gen_reg_1__regIns_N3,
         top_AND_M30_U1_gen_reg_2__regIns_n2,
         top_AND_M30_U1_gen_reg_2__regIns_N3,
         top_AND_M30_U1_gen_reg_3__regIns_n2,
         top_AND_M30_U1_gen_reg_3__regIns_N3,
         top_AND_M30_U1_gen_reg_4__regIns_n2,
         top_AND_M30_U1_gen_reg_4__regIns_N3,
         top_AND_M30_U1_gen_reg_5__regIns_n2,
         top_AND_M30_U1_gen_reg_5__regIns_N3,
         top_AND_M30_U1_gen_reg_6__regIns_n2,
         top_AND_M30_U1_gen_reg_6__regIns_N3,
         top_AND_M30_U1_gen_reg_7__regIns_n2,
         top_AND_M30_U1_gen_reg_7__regIns_N3,
         top_AND_M30_U1_OperationInst_andInst0_n3,
         top_AND_M30_U1_OperationInst_andInst1_n3,
         top_AND_M30_U1_OperationInst_andInst2_n3,
         top_AND_M30_U1_OperationInst_andInst3_n3,
         top_AND_M30_U1_OperationInst_orInst1_n6,
         top_AND_M30_U1_OperationInst_orInst1_n5,
         top_AND_M30_U1_OperationInst_andInst4_n3,
         top_AND_M30_U1_OperationInst_andInst5_n3,
         top_AND_M30_U1_OperationInst_andInst6_n3,
         top_AND_M30_U1_OperationInst_andInst7_n3,
         top_AND_M30_U1_OperationInst_orInst2_n6,
         top_AND_M30_U1_OperationInst_orInst2_n5,
         top_AND_M31_U1_nonlinearInst_n64, top_AND_M31_U1_nonlinearInst_n63,
         top_AND_M31_U1_nonlinearInst_n62, top_AND_M31_U1_nonlinearInst_n61,
         top_AND_M31_U1_nonlinearInst_n60, top_AND_M31_U1_nonlinearInst_n59,
         top_AND_M31_U1_nonlinearInst_n58, top_AND_M31_U1_nonlinearInst_n57,
         top_AND_M31_U1_nonlinearInst_n56, top_AND_M31_U1_nonlinearInst_n55,
         top_AND_M31_U1_nonlinearInst_n54, top_AND_M31_U1_nonlinearInst_n53,
         top_AND_M31_U1_nonlinearInst_n52, top_AND_M31_U1_nonlinearInst_n51,
         top_AND_M31_U1_nonlinearInst_n50, top_AND_M31_U1_nonlinearInst_n49,
         top_AND_M31_U1_nonlinearInst_n48, top_AND_M31_U1_nonlinearInst_n47,
         top_AND_M31_U1_gen_reg_0__regIns_n2,
         top_AND_M31_U1_gen_reg_0__regIns_N3,
         top_AND_M31_U1_gen_reg_1__regIns_n2,
         top_AND_M31_U1_gen_reg_1__regIns_N3,
         top_AND_M31_U1_gen_reg_2__regIns_n2,
         top_AND_M31_U1_gen_reg_2__regIns_N3,
         top_AND_M31_U1_gen_reg_3__regIns_n2,
         top_AND_M31_U1_gen_reg_3__regIns_N3,
         top_AND_M31_U1_gen_reg_4__regIns_n2,
         top_AND_M31_U1_gen_reg_4__regIns_N3,
         top_AND_M31_U1_gen_reg_5__regIns_n2,
         top_AND_M31_U1_gen_reg_5__regIns_N3,
         top_AND_M31_U1_gen_reg_6__regIns_n2,
         top_AND_M31_U1_gen_reg_6__regIns_N3,
         top_AND_M31_U1_gen_reg_7__regIns_n2,
         top_AND_M31_U1_gen_reg_7__regIns_N3,
         top_AND_M31_U1_OperationInst_andInst0_n3,
         top_AND_M31_U1_OperationInst_andInst1_n3,
         top_AND_M31_U1_OperationInst_andInst2_n3,
         top_AND_M31_U1_OperationInst_andInst3_n3,
         top_AND_M31_U1_OperationInst_orInst1_n6,
         top_AND_M31_U1_OperationInst_orInst1_n5,
         top_AND_M31_U1_OperationInst_andInst4_n3,
         top_AND_M31_U1_OperationInst_andInst5_n3,
         top_AND_M31_U1_OperationInst_andInst6_n3,
         top_AND_M31_U1_OperationInst_andInst7_n3,
         top_AND_M31_U1_OperationInst_orInst2_n6,
         top_AND_M31_U1_OperationInst_orInst2_n5,
         top_AND_M32_U1_nonlinearInst_n64, top_AND_M32_U1_nonlinearInst_n63,
         top_AND_M32_U1_nonlinearInst_n62, top_AND_M32_U1_nonlinearInst_n61,
         top_AND_M32_U1_nonlinearInst_n60, top_AND_M32_U1_nonlinearInst_n59,
         top_AND_M32_U1_nonlinearInst_n58, top_AND_M32_U1_nonlinearInst_n57,
         top_AND_M32_U1_nonlinearInst_n56, top_AND_M32_U1_nonlinearInst_n55,
         top_AND_M32_U1_nonlinearInst_n54, top_AND_M32_U1_nonlinearInst_n53,
         top_AND_M32_U1_nonlinearInst_n52, top_AND_M32_U1_nonlinearInst_n51,
         top_AND_M32_U1_nonlinearInst_n50, top_AND_M32_U1_nonlinearInst_n49,
         top_AND_M32_U1_nonlinearInst_n48, top_AND_M32_U1_nonlinearInst_n47,
         top_AND_M32_U1_gen_reg_0__regIns_n2,
         top_AND_M32_U1_gen_reg_0__regIns_N3,
         top_AND_M32_U1_gen_reg_1__regIns_n2,
         top_AND_M32_U1_gen_reg_1__regIns_N3,
         top_AND_M32_U1_gen_reg_2__regIns_n2,
         top_AND_M32_U1_gen_reg_2__regIns_N3,
         top_AND_M32_U1_gen_reg_3__regIns_n2,
         top_AND_M32_U1_gen_reg_3__regIns_N3,
         top_AND_M32_U1_gen_reg_4__regIns_n2,
         top_AND_M32_U1_gen_reg_4__regIns_N3,
         top_AND_M32_U1_gen_reg_5__regIns_n2,
         top_AND_M32_U1_gen_reg_5__regIns_N3,
         top_AND_M32_U1_gen_reg_6__regIns_n2,
         top_AND_M32_U1_gen_reg_6__regIns_N3,
         top_AND_M32_U1_gen_reg_7__regIns_n2,
         top_AND_M32_U1_gen_reg_7__regIns_N3,
         top_AND_M32_U1_OperationInst_andInst0_n3,
         top_AND_M32_U1_OperationInst_andInst1_n3,
         top_AND_M32_U1_OperationInst_andInst2_n3,
         top_AND_M32_U1_OperationInst_andInst3_n3,
         top_AND_M32_U1_OperationInst_orInst1_n6,
         top_AND_M32_U1_OperationInst_orInst1_n5,
         top_AND_M32_U1_OperationInst_andInst4_n3,
         top_AND_M32_U1_OperationInst_andInst5_n3,
         top_AND_M32_U1_OperationInst_andInst6_n3,
         top_AND_M32_U1_OperationInst_andInst7_n3,
         top_AND_M32_U1_OperationInst_orInst2_n6,
         top_AND_M32_U1_OperationInst_orInst2_n5, top_XOR_M33_U1_xorInst_n12,
         top_XOR_M33_U1_xorInst_n11, top_XOR_M33_U1_xorInst_n10,
         top_XOR_M33_U1_xorInst_n9, top_AND_M34_U1_nonlinearInst_n64,
         top_AND_M34_U1_nonlinearInst_n63, top_AND_M34_U1_nonlinearInst_n62,
         top_AND_M34_U1_nonlinearInst_n61, top_AND_M34_U1_nonlinearInst_n60,
         top_AND_M34_U1_nonlinearInst_n59, top_AND_M34_U1_nonlinearInst_n58,
         top_AND_M34_U1_nonlinearInst_n57, top_AND_M34_U1_nonlinearInst_n56,
         top_AND_M34_U1_nonlinearInst_n55, top_AND_M34_U1_nonlinearInst_n54,
         top_AND_M34_U1_nonlinearInst_n53, top_AND_M34_U1_nonlinearInst_n52,
         top_AND_M34_U1_nonlinearInst_n51, top_AND_M34_U1_nonlinearInst_n50,
         top_AND_M34_U1_nonlinearInst_n49, top_AND_M34_U1_nonlinearInst_n48,
         top_AND_M34_U1_nonlinearInst_n47, top_AND_M34_U1_gen_reg_0__regIns_n2,
         top_AND_M34_U1_gen_reg_0__regIns_N3,
         top_AND_M34_U1_gen_reg_1__regIns_n2,
         top_AND_M34_U1_gen_reg_1__regIns_N3,
         top_AND_M34_U1_gen_reg_2__regIns_n2,
         top_AND_M34_U1_gen_reg_2__regIns_N3,
         top_AND_M34_U1_gen_reg_3__regIns_n2,
         top_AND_M34_U1_gen_reg_3__regIns_N3,
         top_AND_M34_U1_gen_reg_4__regIns_n2,
         top_AND_M34_U1_gen_reg_4__regIns_N3,
         top_AND_M34_U1_gen_reg_5__regIns_n2,
         top_AND_M34_U1_gen_reg_5__regIns_N3,
         top_AND_M34_U1_gen_reg_6__regIns_n2,
         top_AND_M34_U1_gen_reg_6__regIns_N3,
         top_AND_M34_U1_gen_reg_7__regIns_n2,
         top_AND_M34_U1_gen_reg_7__regIns_N3,
         top_AND_M34_U1_OperationInst_andInst0_n3,
         top_AND_M34_U1_OperationInst_andInst1_n3,
         top_AND_M34_U1_OperationInst_andInst2_n3,
         top_AND_M34_U1_OperationInst_andInst3_n3,
         top_AND_M34_U1_OperationInst_orInst1_n6,
         top_AND_M34_U1_OperationInst_orInst1_n5,
         top_AND_M34_U1_OperationInst_andInst4_n3,
         top_AND_M34_U1_OperationInst_andInst5_n3,
         top_AND_M34_U1_OperationInst_andInst6_n3,
         top_AND_M34_U1_OperationInst_andInst7_n3,
         top_AND_M34_U1_OperationInst_orInst2_n6,
         top_AND_M34_U1_OperationInst_orInst2_n5,
         top_AND_M35_U1_nonlinearInst_n64, top_AND_M35_U1_nonlinearInst_n63,
         top_AND_M35_U1_nonlinearInst_n62, top_AND_M35_U1_nonlinearInst_n61,
         top_AND_M35_U1_nonlinearInst_n60, top_AND_M35_U1_nonlinearInst_n59,
         top_AND_M35_U1_nonlinearInst_n58, top_AND_M35_U1_nonlinearInst_n57,
         top_AND_M35_U1_nonlinearInst_n56, top_AND_M35_U1_nonlinearInst_n55,
         top_AND_M35_U1_nonlinearInst_n54, top_AND_M35_U1_nonlinearInst_n53,
         top_AND_M35_U1_nonlinearInst_n52, top_AND_M35_U1_nonlinearInst_n51,
         top_AND_M35_U1_nonlinearInst_n50, top_AND_M35_U1_nonlinearInst_n49,
         top_AND_M35_U1_nonlinearInst_n48, top_AND_M35_U1_nonlinearInst_n47,
         top_AND_M35_U1_gen_reg_0__regIns_n2,
         top_AND_M35_U1_gen_reg_0__regIns_N3,
         top_AND_M35_U1_gen_reg_1__regIns_n2,
         top_AND_M35_U1_gen_reg_1__regIns_N3,
         top_AND_M35_U1_gen_reg_2__regIns_n2,
         top_AND_M35_U1_gen_reg_2__regIns_N3,
         top_AND_M35_U1_gen_reg_3__regIns_n2,
         top_AND_M35_U1_gen_reg_3__regIns_N3,
         top_AND_M35_U1_gen_reg_4__regIns_n2,
         top_AND_M35_U1_gen_reg_4__regIns_N3,
         top_AND_M35_U1_gen_reg_5__regIns_n2,
         top_AND_M35_U1_gen_reg_5__regIns_N3,
         top_AND_M35_U1_gen_reg_6__regIns_n2,
         top_AND_M35_U1_gen_reg_6__regIns_N3,
         top_AND_M35_U1_gen_reg_7__regIns_n2,
         top_AND_M35_U1_gen_reg_7__regIns_N3,
         top_AND_M35_U1_OperationInst_andInst0_n3,
         top_AND_M35_U1_OperationInst_andInst1_n3,
         top_AND_M35_U1_OperationInst_andInst2_n3,
         top_AND_M35_U1_OperationInst_andInst3_n3,
         top_AND_M35_U1_OperationInst_orInst1_n6,
         top_AND_M35_U1_OperationInst_orInst1_n5,
         top_AND_M35_U1_OperationInst_andInst4_n3,
         top_AND_M35_U1_OperationInst_andInst5_n3,
         top_AND_M35_U1_OperationInst_andInst6_n3,
         top_AND_M35_U1_OperationInst_andInst7_n3,
         top_AND_M35_U1_OperationInst_orInst2_n6,
         top_AND_M35_U1_OperationInst_orInst2_n5, top_XOR_M36_U1_xorInst_n12,
         top_XOR_M36_U1_xorInst_n11, top_XOR_M36_U1_xorInst_n10,
         top_XOR_M36_U1_xorInst_n9, top_XOR_M37_U1_xorInst_n12,
         top_XOR_M37_U1_xorInst_n11, top_XOR_M37_U1_xorInst_n10,
         top_XOR_M37_U1_xorInst_n9, top_XOR_M38_U1_xorInst_n12,
         top_XOR_M38_U1_xorInst_n11, top_XOR_M38_U1_xorInst_n10,
         top_XOR_M38_U1_xorInst_n9, top_XOR_M39_U1_xorInst_n12,
         top_XOR_M39_U1_xorInst_n11, top_XOR_M39_U1_xorInst_n10,
         top_XOR_M39_U1_xorInst_n9, top_XOR_M40_U1_xorInst_n12,
         top_XOR_M40_U1_xorInst_n11, top_XOR_M40_U1_xorInst_n10,
         top_XOR_M40_U1_xorInst_n9, top_XOR_M41_U1_xorInst_n12,
         top_XOR_M41_U1_xorInst_n11, top_XOR_M41_U1_xorInst_n10,
         top_XOR_M41_U1_xorInst_n9, top_XOR_M42_U1_xorInst_n12,
         top_XOR_M42_U1_xorInst_n11, top_XOR_M42_U1_xorInst_n10,
         top_XOR_M42_U1_xorInst_n9, top_XOR_M43_U1_xorInst_n12,
         top_XOR_M43_U1_xorInst_n11, top_XOR_M43_U1_xorInst_n10,
         top_XOR_M43_U1_xorInst_n9, top_XOR_M44_U1_xorInst_n12,
         top_XOR_M44_U1_xorInst_n11, top_XOR_M44_U1_xorInst_n10,
         top_XOR_M44_U1_xorInst_n9, top_XOR_M45_U1_xorInst_n12,
         top_XOR_M45_U1_xorInst_n11, top_XOR_M45_U1_xorInst_n10,
         top_XOR_M45_U1_xorInst_n9, top_AND_M46_U1_nonlinearInst_n64,
         top_AND_M46_U1_nonlinearInst_n63, top_AND_M46_U1_nonlinearInst_n62,
         top_AND_M46_U1_nonlinearInst_n61, top_AND_M46_U1_nonlinearInst_n60,
         top_AND_M46_U1_nonlinearInst_n59, top_AND_M46_U1_nonlinearInst_n58,
         top_AND_M46_U1_nonlinearInst_n57, top_AND_M46_U1_nonlinearInst_n56,
         top_AND_M46_U1_nonlinearInst_n55, top_AND_M46_U1_nonlinearInst_n54,
         top_AND_M46_U1_nonlinearInst_n53, top_AND_M46_U1_nonlinearInst_n52,
         top_AND_M46_U1_nonlinearInst_n51, top_AND_M46_U1_nonlinearInst_n50,
         top_AND_M46_U1_nonlinearInst_n49, top_AND_M46_U1_nonlinearInst_n48,
         top_AND_M46_U1_nonlinearInst_n47, top_AND_M46_U1_gen_reg_0__regIns_n2,
         top_AND_M46_U1_gen_reg_0__regIns_N3,
         top_AND_M46_U1_gen_reg_1__regIns_n2,
         top_AND_M46_U1_gen_reg_1__regIns_N3,
         top_AND_M46_U1_gen_reg_2__regIns_n2,
         top_AND_M46_U1_gen_reg_2__regIns_N3,
         top_AND_M46_U1_gen_reg_3__regIns_n2,
         top_AND_M46_U1_gen_reg_3__regIns_N3,
         top_AND_M46_U1_gen_reg_4__regIns_n2,
         top_AND_M46_U1_gen_reg_4__regIns_N3,
         top_AND_M46_U1_gen_reg_5__regIns_n2,
         top_AND_M46_U1_gen_reg_5__regIns_N3,
         top_AND_M46_U1_gen_reg_6__regIns_n2,
         top_AND_M46_U1_gen_reg_6__regIns_N3,
         top_AND_M46_U1_gen_reg_7__regIns_n2,
         top_AND_M46_U1_gen_reg_7__regIns_N3,
         top_AND_M46_U1_OperationInst_andInst0_n3,
         top_AND_M46_U1_OperationInst_andInst1_n3,
         top_AND_M46_U1_OperationInst_andInst2_n3,
         top_AND_M46_U1_OperationInst_andInst3_n3,
         top_AND_M46_U1_OperationInst_orInst1_n6,
         top_AND_M46_U1_OperationInst_orInst1_n5,
         top_AND_M46_U1_OperationInst_andInst4_n3,
         top_AND_M46_U1_OperationInst_andInst5_n3,
         top_AND_M46_U1_OperationInst_andInst6_n3,
         top_AND_M46_U1_OperationInst_andInst7_n3,
         top_AND_M46_U1_OperationInst_orInst2_n6,
         top_AND_M46_U1_OperationInst_orInst2_n5,
         top_AND_M47_U1_nonlinearInst_n64, top_AND_M47_U1_nonlinearInst_n63,
         top_AND_M47_U1_nonlinearInst_n62, top_AND_M47_U1_nonlinearInst_n61,
         top_AND_M47_U1_nonlinearInst_n60, top_AND_M47_U1_nonlinearInst_n59,
         top_AND_M47_U1_nonlinearInst_n58, top_AND_M47_U1_nonlinearInst_n57,
         top_AND_M47_U1_nonlinearInst_n56, top_AND_M47_U1_nonlinearInst_n55,
         top_AND_M47_U1_nonlinearInst_n54, top_AND_M47_U1_nonlinearInst_n53,
         top_AND_M47_U1_nonlinearInst_n52, top_AND_M47_U1_nonlinearInst_n51,
         top_AND_M47_U1_nonlinearInst_n50, top_AND_M47_U1_nonlinearInst_n49,
         top_AND_M47_U1_nonlinearInst_n48, top_AND_M47_U1_nonlinearInst_n47,
         top_AND_M47_U1_gen_reg_0__regIns_n2,
         top_AND_M47_U1_gen_reg_0__regIns_N3,
         top_AND_M47_U1_gen_reg_1__regIns_n2,
         top_AND_M47_U1_gen_reg_1__regIns_N3,
         top_AND_M47_U1_gen_reg_2__regIns_n2,
         top_AND_M47_U1_gen_reg_2__regIns_N3,
         top_AND_M47_U1_gen_reg_3__regIns_n2,
         top_AND_M47_U1_gen_reg_3__regIns_N3,
         top_AND_M47_U1_gen_reg_4__regIns_n2,
         top_AND_M47_U1_gen_reg_4__regIns_N3,
         top_AND_M47_U1_gen_reg_5__regIns_n2,
         top_AND_M47_U1_gen_reg_5__regIns_N3,
         top_AND_M47_U1_gen_reg_6__regIns_n2,
         top_AND_M47_U1_gen_reg_6__regIns_N3,
         top_AND_M47_U1_gen_reg_7__regIns_n2,
         top_AND_M47_U1_gen_reg_7__regIns_N3,
         top_AND_M47_U1_OperationInst_andInst0_n3,
         top_AND_M47_U1_OperationInst_andInst1_n3,
         top_AND_M47_U1_OperationInst_andInst2_n3,
         top_AND_M47_U1_OperationInst_andInst3_n3,
         top_AND_M47_U1_OperationInst_orInst1_n6,
         top_AND_M47_U1_OperationInst_orInst1_n5,
         top_AND_M47_U1_OperationInst_andInst4_n3,
         top_AND_M47_U1_OperationInst_andInst5_n3,
         top_AND_M47_U1_OperationInst_andInst6_n3,
         top_AND_M47_U1_OperationInst_andInst7_n3,
         top_AND_M47_U1_OperationInst_orInst2_n6,
         top_AND_M47_U1_OperationInst_orInst2_n5,
         top_AND_M48_U1_nonlinearInst_n64, top_AND_M48_U1_nonlinearInst_n63,
         top_AND_M48_U1_nonlinearInst_n62, top_AND_M48_U1_nonlinearInst_n61,
         top_AND_M48_U1_nonlinearInst_n60, top_AND_M48_U1_nonlinearInst_n59,
         top_AND_M48_U1_nonlinearInst_n58, top_AND_M48_U1_nonlinearInst_n57,
         top_AND_M48_U1_nonlinearInst_n56, top_AND_M48_U1_nonlinearInst_n55,
         top_AND_M48_U1_nonlinearInst_n54, top_AND_M48_U1_nonlinearInst_n53,
         top_AND_M48_U1_nonlinearInst_n52, top_AND_M48_U1_nonlinearInst_n51,
         top_AND_M48_U1_nonlinearInst_n50, top_AND_M48_U1_nonlinearInst_n49,
         top_AND_M48_U1_nonlinearInst_n48, top_AND_M48_U1_nonlinearInst_n47,
         top_AND_M48_U1_gen_reg_0__regIns_n2,
         top_AND_M48_U1_gen_reg_0__regIns_N3,
         top_AND_M48_U1_gen_reg_1__regIns_n2,
         top_AND_M48_U1_gen_reg_1__regIns_N3,
         top_AND_M48_U1_gen_reg_2__regIns_n2,
         top_AND_M48_U1_gen_reg_2__regIns_N3,
         top_AND_M48_U1_gen_reg_3__regIns_n2,
         top_AND_M48_U1_gen_reg_3__regIns_N3,
         top_AND_M48_U1_gen_reg_4__regIns_n2,
         top_AND_M48_U1_gen_reg_4__regIns_N3,
         top_AND_M48_U1_gen_reg_5__regIns_n2,
         top_AND_M48_U1_gen_reg_5__regIns_N3,
         top_AND_M48_U1_gen_reg_6__regIns_n2,
         top_AND_M48_U1_gen_reg_6__regIns_N3,
         top_AND_M48_U1_gen_reg_7__regIns_n2,
         top_AND_M48_U1_gen_reg_7__regIns_N3,
         top_AND_M48_U1_OperationInst_andInst0_n3,
         top_AND_M48_U1_OperationInst_andInst1_n3,
         top_AND_M48_U1_OperationInst_andInst2_n3,
         top_AND_M48_U1_OperationInst_andInst3_n3,
         top_AND_M48_U1_OperationInst_orInst1_n6,
         top_AND_M48_U1_OperationInst_orInst1_n5,
         top_AND_M48_U1_OperationInst_andInst4_n3,
         top_AND_M48_U1_OperationInst_andInst5_n3,
         top_AND_M48_U1_OperationInst_andInst6_n3,
         top_AND_M48_U1_OperationInst_andInst7_n3,
         top_AND_M48_U1_OperationInst_orInst2_n6,
         top_AND_M48_U1_OperationInst_orInst2_n5,
         top_AND_M49_U1_nonlinearInst_n64, top_AND_M49_U1_nonlinearInst_n63,
         top_AND_M49_U1_nonlinearInst_n62, top_AND_M49_U1_nonlinearInst_n61,
         top_AND_M49_U1_nonlinearInst_n60, top_AND_M49_U1_nonlinearInst_n59,
         top_AND_M49_U1_nonlinearInst_n58, top_AND_M49_U1_nonlinearInst_n57,
         top_AND_M49_U1_nonlinearInst_n56, top_AND_M49_U1_nonlinearInst_n55,
         top_AND_M49_U1_nonlinearInst_n54, top_AND_M49_U1_nonlinearInst_n53,
         top_AND_M49_U1_nonlinearInst_n52, top_AND_M49_U1_nonlinearInst_n51,
         top_AND_M49_U1_nonlinearInst_n50, top_AND_M49_U1_nonlinearInst_n49,
         top_AND_M49_U1_nonlinearInst_n48, top_AND_M49_U1_nonlinearInst_n47,
         top_AND_M49_U1_gen_reg_0__regIns_n2,
         top_AND_M49_U1_gen_reg_0__regIns_N3,
         top_AND_M49_U1_gen_reg_1__regIns_n2,
         top_AND_M49_U1_gen_reg_1__regIns_N3,
         top_AND_M49_U1_gen_reg_2__regIns_n2,
         top_AND_M49_U1_gen_reg_2__regIns_N3,
         top_AND_M49_U1_gen_reg_3__regIns_n2,
         top_AND_M49_U1_gen_reg_3__regIns_N3,
         top_AND_M49_U1_gen_reg_4__regIns_n2,
         top_AND_M49_U1_gen_reg_4__regIns_N3,
         top_AND_M49_U1_gen_reg_5__regIns_n2,
         top_AND_M49_U1_gen_reg_5__regIns_N3,
         top_AND_M49_U1_gen_reg_6__regIns_n2,
         top_AND_M49_U1_gen_reg_6__regIns_N3,
         top_AND_M49_U1_gen_reg_7__regIns_n2,
         top_AND_M49_U1_gen_reg_7__regIns_N3,
         top_AND_M49_U1_OperationInst_andInst0_n3,
         top_AND_M49_U1_OperationInst_andInst1_n3,
         top_AND_M49_U1_OperationInst_andInst2_n3,
         top_AND_M49_U1_OperationInst_andInst3_n3,
         top_AND_M49_U1_OperationInst_orInst1_n6,
         top_AND_M49_U1_OperationInst_orInst1_n5,
         top_AND_M49_U1_OperationInst_andInst4_n3,
         top_AND_M49_U1_OperationInst_andInst5_n3,
         top_AND_M49_U1_OperationInst_andInst6_n3,
         top_AND_M49_U1_OperationInst_andInst7_n3,
         top_AND_M49_U1_OperationInst_orInst2_n6,
         top_AND_M49_U1_OperationInst_orInst2_n5,
         top_AND_M50_U1_nonlinearInst_n64, top_AND_M50_U1_nonlinearInst_n63,
         top_AND_M50_U1_nonlinearInst_n62, top_AND_M50_U1_nonlinearInst_n61,
         top_AND_M50_U1_nonlinearInst_n60, top_AND_M50_U1_nonlinearInst_n59,
         top_AND_M50_U1_nonlinearInst_n58, top_AND_M50_U1_nonlinearInst_n57,
         top_AND_M50_U1_nonlinearInst_n56, top_AND_M50_U1_nonlinearInst_n55,
         top_AND_M50_U1_nonlinearInst_n54, top_AND_M50_U1_nonlinearInst_n53,
         top_AND_M50_U1_nonlinearInst_n52, top_AND_M50_U1_nonlinearInst_n51,
         top_AND_M50_U1_nonlinearInst_n50, top_AND_M50_U1_nonlinearInst_n49,
         top_AND_M50_U1_nonlinearInst_n48, top_AND_M50_U1_nonlinearInst_n47,
         top_AND_M50_U1_gen_reg_0__regIns_n2,
         top_AND_M50_U1_gen_reg_0__regIns_N3,
         top_AND_M50_U1_gen_reg_1__regIns_n2,
         top_AND_M50_U1_gen_reg_1__regIns_N3,
         top_AND_M50_U1_gen_reg_2__regIns_n2,
         top_AND_M50_U1_gen_reg_2__regIns_N3,
         top_AND_M50_U1_gen_reg_3__regIns_n2,
         top_AND_M50_U1_gen_reg_3__regIns_N3,
         top_AND_M50_U1_gen_reg_4__regIns_n2,
         top_AND_M50_U1_gen_reg_4__regIns_N3,
         top_AND_M50_U1_gen_reg_5__regIns_n2,
         top_AND_M50_U1_gen_reg_5__regIns_N3,
         top_AND_M50_U1_gen_reg_6__regIns_n2,
         top_AND_M50_U1_gen_reg_6__regIns_N3,
         top_AND_M50_U1_gen_reg_7__regIns_n2,
         top_AND_M50_U1_gen_reg_7__regIns_N3,
         top_AND_M50_U1_OperationInst_andInst0_n3,
         top_AND_M50_U1_OperationInst_andInst1_n3,
         top_AND_M50_U1_OperationInst_andInst2_n3,
         top_AND_M50_U1_OperationInst_andInst3_n3,
         top_AND_M50_U1_OperationInst_orInst1_n6,
         top_AND_M50_U1_OperationInst_orInst1_n5,
         top_AND_M50_U1_OperationInst_andInst4_n3,
         top_AND_M50_U1_OperationInst_andInst5_n3,
         top_AND_M50_U1_OperationInst_andInst6_n3,
         top_AND_M50_U1_OperationInst_andInst7_n3,
         top_AND_M50_U1_OperationInst_orInst2_n6,
         top_AND_M50_U1_OperationInst_orInst2_n5,
         top_AND_M51_U1_nonlinearInst_n64, top_AND_M51_U1_nonlinearInst_n63,
         top_AND_M51_U1_nonlinearInst_n62, top_AND_M51_U1_nonlinearInst_n61,
         top_AND_M51_U1_nonlinearInst_n60, top_AND_M51_U1_nonlinearInst_n59,
         top_AND_M51_U1_nonlinearInst_n58, top_AND_M51_U1_nonlinearInst_n57,
         top_AND_M51_U1_nonlinearInst_n56, top_AND_M51_U1_nonlinearInst_n55,
         top_AND_M51_U1_nonlinearInst_n54, top_AND_M51_U1_nonlinearInst_n53,
         top_AND_M51_U1_nonlinearInst_n52, top_AND_M51_U1_nonlinearInst_n51,
         top_AND_M51_U1_nonlinearInst_n50, top_AND_M51_U1_nonlinearInst_n49,
         top_AND_M51_U1_nonlinearInst_n48, top_AND_M51_U1_nonlinearInst_n47,
         top_AND_M51_U1_gen_reg_0__regIns_n2,
         top_AND_M51_U1_gen_reg_0__regIns_N3,
         top_AND_M51_U1_gen_reg_1__regIns_n2,
         top_AND_M51_U1_gen_reg_1__regIns_N3,
         top_AND_M51_U1_gen_reg_2__regIns_n2,
         top_AND_M51_U1_gen_reg_2__regIns_N3,
         top_AND_M51_U1_gen_reg_3__regIns_n2,
         top_AND_M51_U1_gen_reg_3__regIns_N3,
         top_AND_M51_U1_gen_reg_4__regIns_n2,
         top_AND_M51_U1_gen_reg_4__regIns_N3,
         top_AND_M51_U1_gen_reg_5__regIns_n2,
         top_AND_M51_U1_gen_reg_5__regIns_N3,
         top_AND_M51_U1_gen_reg_6__regIns_n2,
         top_AND_M51_U1_gen_reg_6__regIns_N3,
         top_AND_M51_U1_gen_reg_7__regIns_n2,
         top_AND_M51_U1_gen_reg_7__regIns_N3,
         top_AND_M51_U1_OperationInst_andInst0_n3,
         top_AND_M51_U1_OperationInst_andInst1_n3,
         top_AND_M51_U1_OperationInst_andInst2_n3,
         top_AND_M51_U1_OperationInst_andInst3_n3,
         top_AND_M51_U1_OperationInst_orInst1_n6,
         top_AND_M51_U1_OperationInst_orInst1_n5,
         top_AND_M51_U1_OperationInst_andInst4_n3,
         top_AND_M51_U1_OperationInst_andInst5_n3,
         top_AND_M51_U1_OperationInst_andInst6_n3,
         top_AND_M51_U1_OperationInst_andInst7_n3,
         top_AND_M51_U1_OperationInst_orInst2_n6,
         top_AND_M51_U1_OperationInst_orInst2_n5,
         top_AND_M52_U1_nonlinearInst_n64, top_AND_M52_U1_nonlinearInst_n63,
         top_AND_M52_U1_nonlinearInst_n62, top_AND_M52_U1_nonlinearInst_n61,
         top_AND_M52_U1_nonlinearInst_n60, top_AND_M52_U1_nonlinearInst_n59,
         top_AND_M52_U1_nonlinearInst_n58, top_AND_M52_U1_nonlinearInst_n57,
         top_AND_M52_U1_nonlinearInst_n56, top_AND_M52_U1_nonlinearInst_n55,
         top_AND_M52_U1_nonlinearInst_n54, top_AND_M52_U1_nonlinearInst_n53,
         top_AND_M52_U1_nonlinearInst_n52, top_AND_M52_U1_nonlinearInst_n51,
         top_AND_M52_U1_nonlinearInst_n50, top_AND_M52_U1_nonlinearInst_n49,
         top_AND_M52_U1_nonlinearInst_n48, top_AND_M52_U1_nonlinearInst_n47,
         top_AND_M52_U1_gen_reg_0__regIns_n2,
         top_AND_M52_U1_gen_reg_0__regIns_N3,
         top_AND_M52_U1_gen_reg_1__regIns_n2,
         top_AND_M52_U1_gen_reg_1__regIns_N3,
         top_AND_M52_U1_gen_reg_2__regIns_n2,
         top_AND_M52_U1_gen_reg_2__regIns_N3,
         top_AND_M52_U1_gen_reg_3__regIns_n2,
         top_AND_M52_U1_gen_reg_3__regIns_N3,
         top_AND_M52_U1_gen_reg_4__regIns_n2,
         top_AND_M52_U1_gen_reg_4__regIns_N3,
         top_AND_M52_U1_gen_reg_5__regIns_n2,
         top_AND_M52_U1_gen_reg_5__regIns_N3,
         top_AND_M52_U1_gen_reg_6__regIns_n2,
         top_AND_M52_U1_gen_reg_6__regIns_N3,
         top_AND_M52_U1_gen_reg_7__regIns_n2,
         top_AND_M52_U1_gen_reg_7__regIns_N3,
         top_AND_M52_U1_OperationInst_andInst0_n3,
         top_AND_M52_U1_OperationInst_andInst1_n3,
         top_AND_M52_U1_OperationInst_andInst2_n3,
         top_AND_M52_U1_OperationInst_andInst3_n3,
         top_AND_M52_U1_OperationInst_orInst1_n6,
         top_AND_M52_U1_OperationInst_orInst1_n5,
         top_AND_M52_U1_OperationInst_andInst4_n3,
         top_AND_M52_U1_OperationInst_andInst5_n3,
         top_AND_M52_U1_OperationInst_andInst6_n3,
         top_AND_M52_U1_OperationInst_andInst7_n3,
         top_AND_M52_U1_OperationInst_orInst2_n6,
         top_AND_M52_U1_OperationInst_orInst2_n5,
         top_AND_M53_U1_nonlinearInst_n64, top_AND_M53_U1_nonlinearInst_n63,
         top_AND_M53_U1_nonlinearInst_n62, top_AND_M53_U1_nonlinearInst_n61,
         top_AND_M53_U1_nonlinearInst_n60, top_AND_M53_U1_nonlinearInst_n59,
         top_AND_M53_U1_nonlinearInst_n58, top_AND_M53_U1_nonlinearInst_n57,
         top_AND_M53_U1_nonlinearInst_n56, top_AND_M53_U1_nonlinearInst_n55,
         top_AND_M53_U1_nonlinearInst_n54, top_AND_M53_U1_nonlinearInst_n53,
         top_AND_M53_U1_nonlinearInst_n52, top_AND_M53_U1_nonlinearInst_n51,
         top_AND_M53_U1_nonlinearInst_n50, top_AND_M53_U1_nonlinearInst_n49,
         top_AND_M53_U1_nonlinearInst_n48, top_AND_M53_U1_nonlinearInst_n47,
         top_AND_M53_U1_gen_reg_0__regIns_n2,
         top_AND_M53_U1_gen_reg_0__regIns_N3,
         top_AND_M53_U1_gen_reg_1__regIns_n2,
         top_AND_M53_U1_gen_reg_1__regIns_N3,
         top_AND_M53_U1_gen_reg_2__regIns_n2,
         top_AND_M53_U1_gen_reg_2__regIns_N3,
         top_AND_M53_U1_gen_reg_3__regIns_n2,
         top_AND_M53_U1_gen_reg_3__regIns_N3,
         top_AND_M53_U1_gen_reg_4__regIns_n2,
         top_AND_M53_U1_gen_reg_4__regIns_N3,
         top_AND_M53_U1_gen_reg_5__regIns_n2,
         top_AND_M53_U1_gen_reg_5__regIns_N3,
         top_AND_M53_U1_gen_reg_6__regIns_n2,
         top_AND_M53_U1_gen_reg_6__regIns_N3,
         top_AND_M53_U1_gen_reg_7__regIns_n2,
         top_AND_M53_U1_gen_reg_7__regIns_N3,
         top_AND_M53_U1_OperationInst_andInst0_n3,
         top_AND_M53_U1_OperationInst_andInst1_n3,
         top_AND_M53_U1_OperationInst_andInst2_n3,
         top_AND_M53_U1_OperationInst_andInst3_n3,
         top_AND_M53_U1_OperationInst_orInst1_n6,
         top_AND_M53_U1_OperationInst_orInst1_n5,
         top_AND_M53_U1_OperationInst_andInst4_n3,
         top_AND_M53_U1_OperationInst_andInst5_n3,
         top_AND_M53_U1_OperationInst_andInst6_n3,
         top_AND_M53_U1_OperationInst_andInst7_n3,
         top_AND_M53_U1_OperationInst_orInst2_n6,
         top_AND_M53_U1_OperationInst_orInst2_n5,
         top_AND_M54_U1_nonlinearInst_n64, top_AND_M54_U1_nonlinearInst_n63,
         top_AND_M54_U1_nonlinearInst_n62, top_AND_M54_U1_nonlinearInst_n61,
         top_AND_M54_U1_nonlinearInst_n60, top_AND_M54_U1_nonlinearInst_n59,
         top_AND_M54_U1_nonlinearInst_n58, top_AND_M54_U1_nonlinearInst_n57,
         top_AND_M54_U1_nonlinearInst_n56, top_AND_M54_U1_nonlinearInst_n55,
         top_AND_M54_U1_nonlinearInst_n54, top_AND_M54_U1_nonlinearInst_n53,
         top_AND_M54_U1_nonlinearInst_n52, top_AND_M54_U1_nonlinearInst_n51,
         top_AND_M54_U1_nonlinearInst_n50, top_AND_M54_U1_nonlinearInst_n49,
         top_AND_M54_U1_nonlinearInst_n48, top_AND_M54_U1_nonlinearInst_n47,
         top_AND_M54_U1_gen_reg_0__regIns_n2,
         top_AND_M54_U1_gen_reg_0__regIns_N3,
         top_AND_M54_U1_gen_reg_1__regIns_n2,
         top_AND_M54_U1_gen_reg_1__regIns_N3,
         top_AND_M54_U1_gen_reg_2__regIns_n2,
         top_AND_M54_U1_gen_reg_2__regIns_N3,
         top_AND_M54_U1_gen_reg_3__regIns_n2,
         top_AND_M54_U1_gen_reg_3__regIns_N3,
         top_AND_M54_U1_gen_reg_4__regIns_n2,
         top_AND_M54_U1_gen_reg_4__regIns_N3,
         top_AND_M54_U1_gen_reg_5__regIns_n2,
         top_AND_M54_U1_gen_reg_5__regIns_N3,
         top_AND_M54_U1_gen_reg_6__regIns_n2,
         top_AND_M54_U1_gen_reg_6__regIns_N3,
         top_AND_M54_U1_gen_reg_7__regIns_n2,
         top_AND_M54_U1_gen_reg_7__regIns_N3,
         top_AND_M54_U1_OperationInst_andInst0_n3,
         top_AND_M54_U1_OperationInst_andInst1_n3,
         top_AND_M54_U1_OperationInst_andInst2_n3,
         top_AND_M54_U1_OperationInst_andInst3_n3,
         top_AND_M54_U1_OperationInst_orInst1_n6,
         top_AND_M54_U1_OperationInst_orInst1_n5,
         top_AND_M54_U1_OperationInst_andInst4_n3,
         top_AND_M54_U1_OperationInst_andInst5_n3,
         top_AND_M54_U1_OperationInst_andInst6_n3,
         top_AND_M54_U1_OperationInst_andInst7_n3,
         top_AND_M54_U1_OperationInst_orInst2_n6,
         top_AND_M54_U1_OperationInst_orInst2_n5,
         top_AND_M55_U1_nonlinearInst_n64, top_AND_M55_U1_nonlinearInst_n63,
         top_AND_M55_U1_nonlinearInst_n62, top_AND_M55_U1_nonlinearInst_n61,
         top_AND_M55_U1_nonlinearInst_n60, top_AND_M55_U1_nonlinearInst_n59,
         top_AND_M55_U1_nonlinearInst_n58, top_AND_M55_U1_nonlinearInst_n57,
         top_AND_M55_U1_nonlinearInst_n56, top_AND_M55_U1_nonlinearInst_n55,
         top_AND_M55_U1_nonlinearInst_n54, top_AND_M55_U1_nonlinearInst_n53,
         top_AND_M55_U1_nonlinearInst_n52, top_AND_M55_U1_nonlinearInst_n51,
         top_AND_M55_U1_nonlinearInst_n50, top_AND_M55_U1_nonlinearInst_n49,
         top_AND_M55_U1_nonlinearInst_n48, top_AND_M55_U1_nonlinearInst_n47,
         top_AND_M55_U1_gen_reg_0__regIns_n2,
         top_AND_M55_U1_gen_reg_0__regIns_N3,
         top_AND_M55_U1_gen_reg_1__regIns_n2,
         top_AND_M55_U1_gen_reg_1__regIns_N3,
         top_AND_M55_U1_gen_reg_2__regIns_n2,
         top_AND_M55_U1_gen_reg_2__regIns_N3,
         top_AND_M55_U1_gen_reg_3__regIns_n2,
         top_AND_M55_U1_gen_reg_3__regIns_N3,
         top_AND_M55_U1_gen_reg_4__regIns_n2,
         top_AND_M55_U1_gen_reg_4__regIns_N3,
         top_AND_M55_U1_gen_reg_5__regIns_n2,
         top_AND_M55_U1_gen_reg_5__regIns_N3,
         top_AND_M55_U1_gen_reg_6__regIns_n2,
         top_AND_M55_U1_gen_reg_6__regIns_N3,
         top_AND_M55_U1_gen_reg_7__regIns_n2,
         top_AND_M55_U1_gen_reg_7__regIns_N3,
         top_AND_M55_U1_OperationInst_andInst0_n3,
         top_AND_M55_U1_OperationInst_andInst1_n3,
         top_AND_M55_U1_OperationInst_andInst2_n3,
         top_AND_M55_U1_OperationInst_andInst3_n3,
         top_AND_M55_U1_OperationInst_orInst1_n6,
         top_AND_M55_U1_OperationInst_orInst1_n5,
         top_AND_M55_U1_OperationInst_andInst4_n3,
         top_AND_M55_U1_OperationInst_andInst5_n3,
         top_AND_M55_U1_OperationInst_andInst6_n3,
         top_AND_M55_U1_OperationInst_andInst7_n3,
         top_AND_M55_U1_OperationInst_orInst2_n6,
         top_AND_M55_U1_OperationInst_orInst2_n5,
         top_AND_M56_U1_nonlinearInst_n64, top_AND_M56_U1_nonlinearInst_n63,
         top_AND_M56_U1_nonlinearInst_n62, top_AND_M56_U1_nonlinearInst_n61,
         top_AND_M56_U1_nonlinearInst_n60, top_AND_M56_U1_nonlinearInst_n59,
         top_AND_M56_U1_nonlinearInst_n58, top_AND_M56_U1_nonlinearInst_n57,
         top_AND_M56_U1_nonlinearInst_n56, top_AND_M56_U1_nonlinearInst_n55,
         top_AND_M56_U1_nonlinearInst_n54, top_AND_M56_U1_nonlinearInst_n53,
         top_AND_M56_U1_nonlinearInst_n52, top_AND_M56_U1_nonlinearInst_n51,
         top_AND_M56_U1_nonlinearInst_n50, top_AND_M56_U1_nonlinearInst_n49,
         top_AND_M56_U1_nonlinearInst_n48, top_AND_M56_U1_nonlinearInst_n47,
         top_AND_M56_U1_gen_reg_0__regIns_n2,
         top_AND_M56_U1_gen_reg_0__regIns_N3,
         top_AND_M56_U1_gen_reg_1__regIns_n2,
         top_AND_M56_U1_gen_reg_1__regIns_N3,
         top_AND_M56_U1_gen_reg_2__regIns_n2,
         top_AND_M56_U1_gen_reg_2__regIns_N3,
         top_AND_M56_U1_gen_reg_3__regIns_n2,
         top_AND_M56_U1_gen_reg_3__regIns_N3,
         top_AND_M56_U1_gen_reg_4__regIns_n2,
         top_AND_M56_U1_gen_reg_4__regIns_N3,
         top_AND_M56_U1_gen_reg_5__regIns_n2,
         top_AND_M56_U1_gen_reg_5__regIns_N3,
         top_AND_M56_U1_gen_reg_6__regIns_n2,
         top_AND_M56_U1_gen_reg_6__regIns_N3,
         top_AND_M56_U1_gen_reg_7__regIns_n2,
         top_AND_M56_U1_gen_reg_7__regIns_N3,
         top_AND_M56_U1_OperationInst_andInst0_n3,
         top_AND_M56_U1_OperationInst_andInst1_n3,
         top_AND_M56_U1_OperationInst_andInst2_n3,
         top_AND_M56_U1_OperationInst_andInst3_n3,
         top_AND_M56_U1_OperationInst_orInst1_n6,
         top_AND_M56_U1_OperationInst_orInst1_n5,
         top_AND_M56_U1_OperationInst_andInst4_n3,
         top_AND_M56_U1_OperationInst_andInst5_n3,
         top_AND_M56_U1_OperationInst_andInst6_n3,
         top_AND_M56_U1_OperationInst_andInst7_n3,
         top_AND_M56_U1_OperationInst_orInst2_n6,
         top_AND_M56_U1_OperationInst_orInst2_n5,
         top_AND_M57_U1_nonlinearInst_n64, top_AND_M57_U1_nonlinearInst_n63,
         top_AND_M57_U1_nonlinearInst_n62, top_AND_M57_U1_nonlinearInst_n61,
         top_AND_M57_U1_nonlinearInst_n60, top_AND_M57_U1_nonlinearInst_n59,
         top_AND_M57_U1_nonlinearInst_n58, top_AND_M57_U1_nonlinearInst_n57,
         top_AND_M57_U1_nonlinearInst_n56, top_AND_M57_U1_nonlinearInst_n55,
         top_AND_M57_U1_nonlinearInst_n54, top_AND_M57_U1_nonlinearInst_n53,
         top_AND_M57_U1_nonlinearInst_n52, top_AND_M57_U1_nonlinearInst_n51,
         top_AND_M57_U1_nonlinearInst_n50, top_AND_M57_U1_nonlinearInst_n49,
         top_AND_M57_U1_nonlinearInst_n48, top_AND_M57_U1_nonlinearInst_n47,
         top_AND_M57_U1_gen_reg_0__regIns_n2,
         top_AND_M57_U1_gen_reg_0__regIns_N3,
         top_AND_M57_U1_gen_reg_1__regIns_n2,
         top_AND_M57_U1_gen_reg_1__regIns_N3,
         top_AND_M57_U1_gen_reg_2__regIns_n2,
         top_AND_M57_U1_gen_reg_2__regIns_N3,
         top_AND_M57_U1_gen_reg_3__regIns_n2,
         top_AND_M57_U1_gen_reg_3__regIns_N3,
         top_AND_M57_U1_gen_reg_4__regIns_n2,
         top_AND_M57_U1_gen_reg_4__regIns_N3,
         top_AND_M57_U1_gen_reg_5__regIns_n2,
         top_AND_M57_U1_gen_reg_5__regIns_N3,
         top_AND_M57_U1_gen_reg_6__regIns_n2,
         top_AND_M57_U1_gen_reg_6__regIns_N3,
         top_AND_M57_U1_gen_reg_7__regIns_n2,
         top_AND_M57_U1_gen_reg_7__regIns_N3,
         top_AND_M57_U1_OperationInst_andInst0_n3,
         top_AND_M57_U1_OperationInst_andInst1_n3,
         top_AND_M57_U1_OperationInst_andInst2_n3,
         top_AND_M57_U1_OperationInst_andInst3_n3,
         top_AND_M57_U1_OperationInst_orInst1_n6,
         top_AND_M57_U1_OperationInst_orInst1_n5,
         top_AND_M57_U1_OperationInst_andInst4_n3,
         top_AND_M57_U1_OperationInst_andInst5_n3,
         top_AND_M57_U1_OperationInst_andInst6_n3,
         top_AND_M57_U1_OperationInst_andInst7_n3,
         top_AND_M57_U1_OperationInst_orInst2_n6,
         top_AND_M57_U1_OperationInst_orInst2_n5,
         top_AND_M58_U1_nonlinearInst_n64, top_AND_M58_U1_nonlinearInst_n63,
         top_AND_M58_U1_nonlinearInst_n62, top_AND_M58_U1_nonlinearInst_n61,
         top_AND_M58_U1_nonlinearInst_n60, top_AND_M58_U1_nonlinearInst_n59,
         top_AND_M58_U1_nonlinearInst_n58, top_AND_M58_U1_nonlinearInst_n57,
         top_AND_M58_U1_nonlinearInst_n56, top_AND_M58_U1_nonlinearInst_n55,
         top_AND_M58_U1_nonlinearInst_n54, top_AND_M58_U1_nonlinearInst_n53,
         top_AND_M58_U1_nonlinearInst_n52, top_AND_M58_U1_nonlinearInst_n51,
         top_AND_M58_U1_nonlinearInst_n50, top_AND_M58_U1_nonlinearInst_n49,
         top_AND_M58_U1_nonlinearInst_n48, top_AND_M58_U1_nonlinearInst_n47,
         top_AND_M58_U1_gen_reg_0__regIns_n2,
         top_AND_M58_U1_gen_reg_0__regIns_N3,
         top_AND_M58_U1_gen_reg_1__regIns_n2,
         top_AND_M58_U1_gen_reg_1__regIns_N3,
         top_AND_M58_U1_gen_reg_2__regIns_n2,
         top_AND_M58_U1_gen_reg_2__regIns_N3,
         top_AND_M58_U1_gen_reg_3__regIns_n2,
         top_AND_M58_U1_gen_reg_3__regIns_N3,
         top_AND_M58_U1_gen_reg_4__regIns_n2,
         top_AND_M58_U1_gen_reg_4__regIns_N3,
         top_AND_M58_U1_gen_reg_5__regIns_n2,
         top_AND_M58_U1_gen_reg_5__regIns_N3,
         top_AND_M58_U1_gen_reg_6__regIns_n2,
         top_AND_M58_U1_gen_reg_6__regIns_N3,
         top_AND_M58_U1_gen_reg_7__regIns_n2,
         top_AND_M58_U1_gen_reg_7__regIns_N3,
         top_AND_M58_U1_OperationInst_andInst0_n3,
         top_AND_M58_U1_OperationInst_andInst1_n3,
         top_AND_M58_U1_OperationInst_andInst2_n3,
         top_AND_M58_U1_OperationInst_andInst3_n3,
         top_AND_M58_U1_OperationInst_orInst1_n6,
         top_AND_M58_U1_OperationInst_orInst1_n5,
         top_AND_M58_U1_OperationInst_andInst4_n3,
         top_AND_M58_U1_OperationInst_andInst5_n3,
         top_AND_M58_U1_OperationInst_andInst6_n3,
         top_AND_M58_U1_OperationInst_andInst7_n3,
         top_AND_M58_U1_OperationInst_orInst2_n6,
         top_AND_M58_U1_OperationInst_orInst2_n5,
         top_AND_M59_U1_nonlinearInst_n64, top_AND_M59_U1_nonlinearInst_n63,
         top_AND_M59_U1_nonlinearInst_n62, top_AND_M59_U1_nonlinearInst_n61,
         top_AND_M59_U1_nonlinearInst_n60, top_AND_M59_U1_nonlinearInst_n59,
         top_AND_M59_U1_nonlinearInst_n58, top_AND_M59_U1_nonlinearInst_n57,
         top_AND_M59_U1_nonlinearInst_n56, top_AND_M59_U1_nonlinearInst_n55,
         top_AND_M59_U1_nonlinearInst_n54, top_AND_M59_U1_nonlinearInst_n53,
         top_AND_M59_U1_nonlinearInst_n52, top_AND_M59_U1_nonlinearInst_n51,
         top_AND_M59_U1_nonlinearInst_n50, top_AND_M59_U1_nonlinearInst_n49,
         top_AND_M59_U1_nonlinearInst_n48, top_AND_M59_U1_nonlinearInst_n47,
         top_AND_M59_U1_gen_reg_0__regIns_n2,
         top_AND_M59_U1_gen_reg_0__regIns_N3,
         top_AND_M59_U1_gen_reg_1__regIns_n2,
         top_AND_M59_U1_gen_reg_1__regIns_N3,
         top_AND_M59_U1_gen_reg_2__regIns_n2,
         top_AND_M59_U1_gen_reg_2__regIns_N3,
         top_AND_M59_U1_gen_reg_3__regIns_n2,
         top_AND_M59_U1_gen_reg_3__regIns_N3,
         top_AND_M59_U1_gen_reg_4__regIns_n2,
         top_AND_M59_U1_gen_reg_4__regIns_N3,
         top_AND_M59_U1_gen_reg_5__regIns_n2,
         top_AND_M59_U1_gen_reg_5__regIns_N3,
         top_AND_M59_U1_gen_reg_6__regIns_n2,
         top_AND_M59_U1_gen_reg_6__regIns_N3,
         top_AND_M59_U1_gen_reg_7__regIns_n2,
         top_AND_M59_U1_gen_reg_7__regIns_N3,
         top_AND_M59_U1_OperationInst_andInst0_n3,
         top_AND_M59_U1_OperationInst_andInst1_n3,
         top_AND_M59_U1_OperationInst_andInst2_n3,
         top_AND_M59_U1_OperationInst_andInst3_n3,
         top_AND_M59_U1_OperationInst_orInst1_n6,
         top_AND_M59_U1_OperationInst_orInst1_n5,
         top_AND_M59_U1_OperationInst_andInst4_n3,
         top_AND_M59_U1_OperationInst_andInst5_n3,
         top_AND_M59_U1_OperationInst_andInst6_n3,
         top_AND_M59_U1_OperationInst_andInst7_n3,
         top_AND_M59_U1_OperationInst_orInst2_n6,
         top_AND_M59_U1_OperationInst_orInst2_n5,
         top_AND_M60_U1_nonlinearInst_n64, top_AND_M60_U1_nonlinearInst_n63,
         top_AND_M60_U1_nonlinearInst_n62, top_AND_M60_U1_nonlinearInst_n61,
         top_AND_M60_U1_nonlinearInst_n60, top_AND_M60_U1_nonlinearInst_n59,
         top_AND_M60_U1_nonlinearInst_n58, top_AND_M60_U1_nonlinearInst_n57,
         top_AND_M60_U1_nonlinearInst_n56, top_AND_M60_U1_nonlinearInst_n55,
         top_AND_M60_U1_nonlinearInst_n54, top_AND_M60_U1_nonlinearInst_n53,
         top_AND_M60_U1_nonlinearInst_n52, top_AND_M60_U1_nonlinearInst_n51,
         top_AND_M60_U1_nonlinearInst_n50, top_AND_M60_U1_nonlinearInst_n49,
         top_AND_M60_U1_nonlinearInst_n48, top_AND_M60_U1_nonlinearInst_n47,
         top_AND_M60_U1_gen_reg_0__regIns_n2,
         top_AND_M60_U1_gen_reg_0__regIns_N3,
         top_AND_M60_U1_gen_reg_1__regIns_n2,
         top_AND_M60_U1_gen_reg_1__regIns_N3,
         top_AND_M60_U1_gen_reg_2__regIns_n2,
         top_AND_M60_U1_gen_reg_2__regIns_N3,
         top_AND_M60_U1_gen_reg_3__regIns_n2,
         top_AND_M60_U1_gen_reg_3__regIns_N3,
         top_AND_M60_U1_gen_reg_4__regIns_n2,
         top_AND_M60_U1_gen_reg_4__regIns_N3,
         top_AND_M60_U1_gen_reg_5__regIns_n2,
         top_AND_M60_U1_gen_reg_5__regIns_N3,
         top_AND_M60_U1_gen_reg_6__regIns_n2,
         top_AND_M60_U1_gen_reg_6__regIns_N3,
         top_AND_M60_U1_gen_reg_7__regIns_n2,
         top_AND_M60_U1_gen_reg_7__regIns_N3,
         top_AND_M60_U1_OperationInst_andInst0_n3,
         top_AND_M60_U1_OperationInst_andInst1_n3,
         top_AND_M60_U1_OperationInst_andInst2_n3,
         top_AND_M60_U1_OperationInst_andInst3_n3,
         top_AND_M60_U1_OperationInst_orInst1_n6,
         top_AND_M60_U1_OperationInst_orInst1_n5,
         top_AND_M60_U1_OperationInst_andInst4_n3,
         top_AND_M60_U1_OperationInst_andInst5_n3,
         top_AND_M60_U1_OperationInst_andInst6_n3,
         top_AND_M60_U1_OperationInst_andInst7_n3,
         top_AND_M60_U1_OperationInst_orInst2_n6,
         top_AND_M60_U1_OperationInst_orInst2_n5,
         top_AND_M61_U1_nonlinearInst_n64, top_AND_M61_U1_nonlinearInst_n63,
         top_AND_M61_U1_nonlinearInst_n62, top_AND_M61_U1_nonlinearInst_n61,
         top_AND_M61_U1_nonlinearInst_n60, top_AND_M61_U1_nonlinearInst_n59,
         top_AND_M61_U1_nonlinearInst_n58, top_AND_M61_U1_nonlinearInst_n57,
         top_AND_M61_U1_nonlinearInst_n56, top_AND_M61_U1_nonlinearInst_n55,
         top_AND_M61_U1_nonlinearInst_n54, top_AND_M61_U1_nonlinearInst_n53,
         top_AND_M61_U1_nonlinearInst_n52, top_AND_M61_U1_nonlinearInst_n51,
         top_AND_M61_U1_nonlinearInst_n50, top_AND_M61_U1_nonlinearInst_n49,
         top_AND_M61_U1_nonlinearInst_n48, top_AND_M61_U1_nonlinearInst_n47,
         top_AND_M61_U1_gen_reg_0__regIns_n2,
         top_AND_M61_U1_gen_reg_0__regIns_N3,
         top_AND_M61_U1_gen_reg_1__regIns_n2,
         top_AND_M61_U1_gen_reg_1__regIns_N3,
         top_AND_M61_U1_gen_reg_2__regIns_n2,
         top_AND_M61_U1_gen_reg_2__regIns_N3,
         top_AND_M61_U1_gen_reg_3__regIns_n2,
         top_AND_M61_U1_gen_reg_3__regIns_N3,
         top_AND_M61_U1_gen_reg_4__regIns_n2,
         top_AND_M61_U1_gen_reg_4__regIns_N3,
         top_AND_M61_U1_gen_reg_5__regIns_n2,
         top_AND_M61_U1_gen_reg_5__regIns_N3,
         top_AND_M61_U1_gen_reg_6__regIns_n2,
         top_AND_M61_U1_gen_reg_6__regIns_N3,
         top_AND_M61_U1_gen_reg_7__regIns_n2,
         top_AND_M61_U1_gen_reg_7__regIns_N3,
         top_AND_M61_U1_OperationInst_andInst0_n3,
         top_AND_M61_U1_OperationInst_andInst1_n3,
         top_AND_M61_U1_OperationInst_andInst2_n3,
         top_AND_M61_U1_OperationInst_andInst3_n3,
         top_AND_M61_U1_OperationInst_orInst1_n6,
         top_AND_M61_U1_OperationInst_orInst1_n5,
         top_AND_M61_U1_OperationInst_andInst4_n3,
         top_AND_M61_U1_OperationInst_andInst5_n3,
         top_AND_M61_U1_OperationInst_andInst6_n3,
         top_AND_M61_U1_OperationInst_andInst7_n3,
         top_AND_M61_U1_OperationInst_orInst2_n6,
         top_AND_M61_U1_OperationInst_orInst2_n5,
         top_AND_M62_U1_nonlinearInst_n64, top_AND_M62_U1_nonlinearInst_n63,
         top_AND_M62_U1_nonlinearInst_n62, top_AND_M62_U1_nonlinearInst_n61,
         top_AND_M62_U1_nonlinearInst_n60, top_AND_M62_U1_nonlinearInst_n59,
         top_AND_M62_U1_nonlinearInst_n58, top_AND_M62_U1_nonlinearInst_n57,
         top_AND_M62_U1_nonlinearInst_n56, top_AND_M62_U1_nonlinearInst_n55,
         top_AND_M62_U1_nonlinearInst_n54, top_AND_M62_U1_nonlinearInst_n53,
         top_AND_M62_U1_nonlinearInst_n52, top_AND_M62_U1_nonlinearInst_n51,
         top_AND_M62_U1_nonlinearInst_n50, top_AND_M62_U1_nonlinearInst_n49,
         top_AND_M62_U1_nonlinearInst_n48, top_AND_M62_U1_nonlinearInst_n47,
         top_AND_M62_U1_gen_reg_0__regIns_n2,
         top_AND_M62_U1_gen_reg_0__regIns_N3,
         top_AND_M62_U1_gen_reg_1__regIns_n2,
         top_AND_M62_U1_gen_reg_1__regIns_N3,
         top_AND_M62_U1_gen_reg_2__regIns_n2,
         top_AND_M62_U1_gen_reg_2__regIns_N3,
         top_AND_M62_U1_gen_reg_3__regIns_n2,
         top_AND_M62_U1_gen_reg_3__regIns_N3,
         top_AND_M62_U1_gen_reg_4__regIns_n2,
         top_AND_M62_U1_gen_reg_4__regIns_N3,
         top_AND_M62_U1_gen_reg_5__regIns_n2,
         top_AND_M62_U1_gen_reg_5__regIns_N3,
         top_AND_M62_U1_gen_reg_6__regIns_n2,
         top_AND_M62_U1_gen_reg_6__regIns_N3,
         top_AND_M62_U1_gen_reg_7__regIns_n2,
         top_AND_M62_U1_gen_reg_7__regIns_N3,
         top_AND_M62_U1_OperationInst_andInst0_n3,
         top_AND_M62_U1_OperationInst_andInst1_n3,
         top_AND_M62_U1_OperationInst_andInst2_n3,
         top_AND_M62_U1_OperationInst_andInst3_n3,
         top_AND_M62_U1_OperationInst_orInst1_n6,
         top_AND_M62_U1_OperationInst_orInst1_n5,
         top_AND_M62_U1_OperationInst_andInst4_n3,
         top_AND_M62_U1_OperationInst_andInst5_n3,
         top_AND_M62_U1_OperationInst_andInst6_n3,
         top_AND_M62_U1_OperationInst_andInst7_n3,
         top_AND_M62_U1_OperationInst_orInst2_n6,
         top_AND_M62_U1_OperationInst_orInst2_n5,
         top_AND_M63_U1_nonlinearInst_n64, top_AND_M63_U1_nonlinearInst_n63,
         top_AND_M63_U1_nonlinearInst_n62, top_AND_M63_U1_nonlinearInst_n61,
         top_AND_M63_U1_nonlinearInst_n60, top_AND_M63_U1_nonlinearInst_n59,
         top_AND_M63_U1_nonlinearInst_n58, top_AND_M63_U1_nonlinearInst_n57,
         top_AND_M63_U1_nonlinearInst_n56, top_AND_M63_U1_nonlinearInst_n55,
         top_AND_M63_U1_nonlinearInst_n54, top_AND_M63_U1_nonlinearInst_n53,
         top_AND_M63_U1_nonlinearInst_n52, top_AND_M63_U1_nonlinearInst_n51,
         top_AND_M63_U1_nonlinearInst_n50, top_AND_M63_U1_nonlinearInst_n49,
         top_AND_M63_U1_nonlinearInst_n48, top_AND_M63_U1_nonlinearInst_n47,
         top_AND_M63_U1_gen_reg_0__regIns_n2,
         top_AND_M63_U1_gen_reg_0__regIns_N3,
         top_AND_M63_U1_gen_reg_1__regIns_n2,
         top_AND_M63_U1_gen_reg_1__regIns_N3,
         top_AND_M63_U1_gen_reg_2__regIns_n2,
         top_AND_M63_U1_gen_reg_2__regIns_N3,
         top_AND_M63_U1_gen_reg_3__regIns_n2,
         top_AND_M63_U1_gen_reg_3__regIns_N3,
         top_AND_M63_U1_gen_reg_4__regIns_n2,
         top_AND_M63_U1_gen_reg_4__regIns_N3,
         top_AND_M63_U1_gen_reg_5__regIns_n2,
         top_AND_M63_U1_gen_reg_5__regIns_N3,
         top_AND_M63_U1_gen_reg_6__regIns_n2,
         top_AND_M63_U1_gen_reg_6__regIns_N3,
         top_AND_M63_U1_gen_reg_7__regIns_n2,
         top_AND_M63_U1_gen_reg_7__regIns_N3,
         top_AND_M63_U1_OperationInst_andInst0_n3,
         top_AND_M63_U1_OperationInst_andInst1_n3,
         top_AND_M63_U1_OperationInst_andInst2_n3,
         top_AND_M63_U1_OperationInst_andInst3_n3,
         top_AND_M63_U1_OperationInst_orInst1_n6,
         top_AND_M63_U1_OperationInst_orInst1_n5,
         top_AND_M63_U1_OperationInst_andInst4_n3,
         top_AND_M63_U1_OperationInst_andInst5_n3,
         top_AND_M63_U1_OperationInst_andInst6_n3,
         top_AND_M63_U1_OperationInst_andInst7_n3,
         top_AND_M63_U1_OperationInst_orInst2_n6,
         top_AND_M63_U1_OperationInst_orInst2_n5, top_XOR_L0_U1_xorInst_n12,
         top_XOR_L0_U1_xorInst_n11, top_XOR_L0_U1_xorInst_n10,
         top_XOR_L0_U1_xorInst_n9, top_XOR_L1_U1_xorInst_n12,
         top_XOR_L1_U1_xorInst_n11, top_XOR_L1_U1_xorInst_n10,
         top_XOR_L1_U1_xorInst_n9, top_XOR_L2_U1_xorInst_n12,
         top_XOR_L2_U1_xorInst_n11, top_XOR_L2_U1_xorInst_n10,
         top_XOR_L2_U1_xorInst_n9, top_XOR_L3_U1_xorInst_n12,
         top_XOR_L3_U1_xorInst_n11, top_XOR_L3_U1_xorInst_n10,
         top_XOR_L3_U1_xorInst_n9, top_XOR_L4_U1_xorInst_n12,
         top_XOR_L4_U1_xorInst_n11, top_XOR_L4_U1_xorInst_n10,
         top_XOR_L4_U1_xorInst_n9, top_XOR_L5_U1_xorInst_n12,
         top_XOR_L5_U1_xorInst_n11, top_XOR_L5_U1_xorInst_n10,
         top_XOR_L5_U1_xorInst_n9, top_XOR_L6_U1_xorInst_n12,
         top_XOR_L6_U1_xorInst_n11, top_XOR_L6_U1_xorInst_n10,
         top_XOR_L6_U1_xorInst_n9, top_XOR_L7_U1_xorInst_n12,
         top_XOR_L7_U1_xorInst_n11, top_XOR_L7_U1_xorInst_n10,
         top_XOR_L7_U1_xorInst_n9, top_XOR_L8_U1_xorInst_n12,
         top_XOR_L8_U1_xorInst_n11, top_XOR_L8_U1_xorInst_n10,
         top_XOR_L8_U1_xorInst_n9, top_XOR_L9_U1_xorInst_n12,
         top_XOR_L9_U1_xorInst_n11, top_XOR_L9_U1_xorInst_n10,
         top_XOR_L9_U1_xorInst_n9, top_XOR_L10_U1_xorInst_n12,
         top_XOR_L10_U1_xorInst_n11, top_XOR_L10_U1_xorInst_n10,
         top_XOR_L10_U1_xorInst_n9, top_XOR_L11_U1_xorInst_n12,
         top_XOR_L11_U1_xorInst_n11, top_XOR_L11_U1_xorInst_n10,
         top_XOR_L11_U1_xorInst_n9, top_XOR_L12_U1_xorInst_n12,
         top_XOR_L12_U1_xorInst_n11, top_XOR_L12_U1_xorInst_n10,
         top_XOR_L12_U1_xorInst_n9, top_XOR_L13_U1_xorInst_n12,
         top_XOR_L13_U1_xorInst_n11, top_XOR_L13_U1_xorInst_n10,
         top_XOR_L13_U1_xorInst_n9, top_XOR_L14_U1_xorInst_n12,
         top_XOR_L14_U1_xorInst_n11, top_XOR_L14_U1_xorInst_n10,
         top_XOR_L14_U1_xorInst_n9, top_XOR_L15_U1_xorInst_n12,
         top_XOR_L15_U1_xorInst_n11, top_XOR_L15_U1_xorInst_n10,
         top_XOR_L15_U1_xorInst_n9, top_XOR_L16_U1_xorInst_n12,
         top_XOR_L16_U1_xorInst_n11, top_XOR_L16_U1_xorInst_n10,
         top_XOR_L16_U1_xorInst_n9, top_XOR_L17_U1_xorInst_n12,
         top_XOR_L17_U1_xorInst_n11, top_XOR_L17_U1_xorInst_n10,
         top_XOR_L17_U1_xorInst_n9, top_XOR_L18_U1_xorInst_n12,
         top_XOR_L18_U1_xorInst_n11, top_XOR_L18_U1_xorInst_n10,
         top_XOR_L18_U1_xorInst_n9, top_XOR_L19_U1_xorInst_n12,
         top_XOR_L19_U1_xorInst_n11, top_XOR_L19_U1_xorInst_n10,
         top_XOR_L19_U1_xorInst_n9, top_XOR_L20_U1_xorInst_n12,
         top_XOR_L20_U1_xorInst_n11, top_XOR_L20_U1_xorInst_n10,
         top_XOR_L20_U1_xorInst_n9, top_XOR_L21_U1_xorInst_n12,
         top_XOR_L21_U1_xorInst_n11, top_XOR_L21_U1_xorInst_n10,
         top_XOR_L21_U1_xorInst_n9, top_XOR_L22_U1_xorInst_n12,
         top_XOR_L22_U1_xorInst_n11, top_XOR_L22_U1_xorInst_n10,
         top_XOR_L22_U1_xorInst_n9, top_XOR_L23_U1_xorInst_n12,
         top_XOR_L23_U1_xorInst_n11, top_XOR_L23_U1_xorInst_n10,
         top_XOR_L23_U1_xorInst_n9, top_XOR_L24_U1_xorInst_n12,
         top_XOR_L24_U1_xorInst_n11, top_XOR_L24_U1_xorInst_n10,
         top_XOR_L24_U1_xorInst_n9, top_XOR_L25_U1_xorInst_n12,
         top_XOR_L25_U1_xorInst_n11, top_XOR_L25_U1_xorInst_n10,
         top_XOR_L25_U1_xorInst_n9, top_XOR_L26_U1_xorInst_n12,
         top_XOR_L26_U1_xorInst_n11, top_XOR_L26_U1_xorInst_n10,
         top_XOR_L26_U1_xorInst_n9, top_XOR_L27_U1_xorInst_n12,
         top_XOR_L27_U1_xorInst_n11, top_XOR_L27_U1_xorInst_n10,
         top_XOR_L27_U1_xorInst_n9, top_XOR_L28_U1_xorInst_n12,
         top_XOR_L28_U1_xorInst_n11, top_XOR_L28_U1_xorInst_n10,
         top_XOR_L28_U1_xorInst_n9, top_XOR_L29_U1_xorInst_n12,
         top_XOR_L29_U1_xorInst_n11, top_XOR_L29_U1_xorInst_n10,
         top_XOR_L29_U1_xorInst_n9, top_XOR_S0_U1_c_2_,
         top_XOR_S0_U1_xorInst_n12, top_XOR_S0_U1_xorInst_n11,
         top_XOR_S0_U1_xorInst_n10, top_XOR_S0_U1_xorInst_n9,
         top_XOR_S1_U1_c_2_, top_XOR_S1_U1_xorInst_n12,
         top_XOR_S1_U1_xorInst_n11, top_XOR_S1_U1_xorInst_n10,
         top_XOR_S1_U1_xorInst_n9, top_XOR_S2_U1_c_2_,
         top_XOR_S2_U1_xorInst_n12, top_XOR_S2_U1_xorInst_n11,
         top_XOR_S2_U1_xorInst_n10, top_XOR_S2_U1_xorInst_n9,
         top_XOR_S3_U1_c_2_, top_XOR_S3_U1_xorInst_n12,
         top_XOR_S3_U1_xorInst_n11, top_XOR_S3_U1_xorInst_n10,
         top_XOR_S3_U1_xorInst_n9, top_XOR_S4_U1_c_2_,
         top_XOR_S4_U1_xorInst_n12, top_XOR_S4_U1_xorInst_n11,
         top_XOR_S4_U1_xorInst_n10, top_XOR_S4_U1_xorInst_n9,
         top_XOR_S5_U1_c_2_, top_XOR_S5_U1_xorInst_n12,
         top_XOR_S5_U1_xorInst_n11, top_XOR_S5_U1_xorInst_n10,
         top_XOR_S5_U1_xorInst_n9, top_XOR_S6_U1_c_2_,
         top_XOR_S6_U1_xorInst_n12, top_XOR_S6_U1_xorInst_n11,
         top_XOR_S6_U1_xorInst_n10, top_XOR_S6_U1_xorInst_n9,
         top_XOR_S7_U1_c_2_, top_XOR_S7_U1_xorInst_n12,
         top_XOR_S7_U1_xorInst_n11, top_XOR_S7_U1_xorInst_n10,
         top_XOR_S7_U1_xorInst_n9;
  wire   [3:0] top_XOR_T1_U1_w;
  wire   [3:0] top_XOR_T2_U1_w;
  wire   [3:0] top_XOR_T3_U1_w;
  wire   [3:0] top_XOR_T4_U1_w;
  wire   [3:0] top_XOR_T5_U1_w;
  wire   [3:0] top_XOR_T6_U1_w;
  wire   [3:0] top_XOR_T7_U1_w;
  wire   [3:0] top_XOR_T8_U1_w;
  wire   [3:0] top_XOR_T9_U1_w;
  wire   [3:0] top_XOR_T10_U1_w;
  wire   [3:0] top_XOR_T11_U1_w;
  wire   [3:0] top_XOR_T12_U1_w;
  wire   [3:0] top_XOR_T13_U1_w;
  wire   [3:0] top_XOR_T14_U1_w;
  wire   [3:0] top_XOR_T15_U1_w;
  wire   [3:0] top_XOR_T16_U1_w;
  wire   [3:0] top_XOR_T17_U1_w;
  wire   [3:0] top_XOR_T18_U1_w;
  wire   [3:0] top_XOR_T19_U1_w;
  wire   [3:0] top_XOR_T20_U1_w;
  wire   [3:0] top_XOR_T21_U1_w;
  wire   [3:0] top_XOR_T22_U1_w;
  wire   [3:0] top_XOR_T23_U1_w;
  wire   [3:0] top_XOR_T24_U1_w;
  wire   [3:0] top_XOR_T25_U1_w;
  wire   [3:0] top_XOR_T26_U1_w;
  wire   [3:0] top_XOR_T27_U1_w;
  wire   [7:0] top_AND_M1_U1_t_reg;
  wire   [7:0] top_AND_M1_U1_t;
  wire   [7:0] top_AND_M1_U1_OperationInst_q;
  wire   [7:0] top_AND_M2_U1_t_reg;
  wire   [7:0] top_AND_M2_U1_t;
  wire   [7:0] top_AND_M2_U1_OperationInst_q;
  wire   [3:0] top_XOR_M3_U1_w;
  wire   [7:0] top_AND_M4_U1_t_reg;
  wire   [7:0] top_AND_M4_U1_t;
  wire   [7:0] top_AND_M4_U1_OperationInst_q;
  wire   [3:0] top_XOR_M5_U1_w;
  wire   [7:0] top_AND_M6_U1_t_reg;
  wire   [7:0] top_AND_M6_U1_t;
  wire   [7:0] top_AND_M6_U1_OperationInst_q;
  wire   [7:0] top_AND_M7_U1_t_reg;
  wire   [7:0] top_AND_M7_U1_t;
  wire   [7:0] top_AND_M7_U1_OperationInst_q;
  wire   [3:0] top_XOR_M8_U1_w;
  wire   [7:0] top_AND_M9_U1_t_reg;
  wire   [7:0] top_AND_M9_U1_t;
  wire   [7:0] top_AND_M9_U1_OperationInst_q;
  wire   [3:0] top_XOR_M10_U1_w;
  wire   [7:0] top_AND_M11_U1_t_reg;
  wire   [7:0] top_AND_M11_U1_t;
  wire   [7:0] top_AND_M11_U1_OperationInst_q;
  wire   [7:0] top_AND_M12_U1_t_reg;
  wire   [7:0] top_AND_M12_U1_t;
  wire   [7:0] top_AND_M12_U1_OperationInst_q;
  wire   [3:0] top_XOR_M13_U1_w;
  wire   [7:0] top_AND_M14_U1_t_reg;
  wire   [7:0] top_AND_M14_U1_t;
  wire   [7:0] top_AND_M14_U1_OperationInst_q;
  wire   [3:0] top_XOR_M15_U1_w;
  wire   [3:0] top_XOR_M16_U1_w;
  wire   [3:0] top_XOR_M17_U1_w;
  wire   [3:0] top_XOR_M18_U1_w;
  wire   [3:0] top_XOR_M19_U1_w;
  wire   [3:0] top_XOR_M20_U1_w;
  wire   [3:0] top_XOR_M21_U1_w;
  wire   [3:0] top_XOR_M22_U1_w;
  wire   [3:0] top_XOR_M23_U1_w;
  wire   [3:0] top_XOR_M24_U1_w;
  wire   [7:0] top_AND_M25_U1_t_reg;
  wire   [7:0] top_AND_M25_U1_t;
  wire   [7:0] top_AND_M25_U1_OperationInst_q;
  wire   [3:0] top_XOR_M26_U1_w;
  wire   [3:0] top_XOR_M27_U1_w;
  wire   [3:0] top_XOR_M28_U1_w;
  wire   [7:0] top_AND_M29_U1_t_reg;
  wire   [7:0] top_AND_M29_U1_t;
  wire   [7:0] top_AND_M29_U1_OperationInst_q;
  wire   [7:0] top_AND_M30_U1_t_reg;
  wire   [7:0] top_AND_M30_U1_t;
  wire   [7:0] top_AND_M30_U1_OperationInst_q;
  wire   [7:0] top_AND_M31_U1_t_reg;
  wire   [7:0] top_AND_M31_U1_t;
  wire   [7:0] top_AND_M31_U1_OperationInst_q;
  wire   [7:0] top_AND_M32_U1_t_reg;
  wire   [7:0] top_AND_M32_U1_t;
  wire   [7:0] top_AND_M32_U1_OperationInst_q;
  wire   [3:0] top_XOR_M33_U1_w;
  wire   [7:0] top_AND_M34_U1_t_reg;
  wire   [7:0] top_AND_M34_U1_t;
  wire   [7:0] top_AND_M34_U1_OperationInst_q;
  wire   [7:0] top_AND_M35_U1_t_reg;
  wire   [7:0] top_AND_M35_U1_t;
  wire   [7:0] top_AND_M35_U1_OperationInst_q;
  wire   [3:0] top_XOR_M36_U1_w;
  wire   [3:0] top_XOR_M37_U1_w;
  wire   [3:0] top_XOR_M38_U1_w;
  wire   [3:0] top_XOR_M39_U1_w;
  wire   [3:0] top_XOR_M40_U1_w;
  wire   [3:0] top_XOR_M41_U1_w;
  wire   [3:0] top_XOR_M42_U1_w;
  wire   [3:0] top_XOR_M43_U1_w;
  wire   [3:0] top_XOR_M44_U1_w;
  wire   [3:0] top_XOR_M45_U1_w;
  wire   [7:0] top_AND_M46_U1_t_reg;
  wire   [7:0] top_AND_M46_U1_t;
  wire   [7:0] top_AND_M46_U1_OperationInst_q;
  wire   [7:0] top_AND_M47_U1_t_reg;
  wire   [7:0] top_AND_M47_U1_t;
  wire   [7:0] top_AND_M47_U1_OperationInst_q;
  wire   [7:0] top_AND_M48_U1_t_reg;
  wire   [7:0] top_AND_M48_U1_t;
  wire   [7:0] top_AND_M48_U1_OperationInst_q;
  wire   [7:0] top_AND_M49_U1_t_reg;
  wire   [7:0] top_AND_M49_U1_t;
  wire   [7:0] top_AND_M49_U1_OperationInst_q;
  wire   [7:0] top_AND_M50_U1_t_reg;
  wire   [7:0] top_AND_M50_U1_t;
  wire   [7:0] top_AND_M50_U1_OperationInst_q;
  wire   [7:0] top_AND_M51_U1_t_reg;
  wire   [7:0] top_AND_M51_U1_t;
  wire   [7:0] top_AND_M51_U1_OperationInst_q;
  wire   [7:0] top_AND_M52_U1_t_reg;
  wire   [7:0] top_AND_M52_U1_t;
  wire   [7:0] top_AND_M52_U1_OperationInst_q;
  wire   [7:0] top_AND_M53_U1_t_reg;
  wire   [7:0] top_AND_M53_U1_t;
  wire   [7:0] top_AND_M53_U1_OperationInst_q;
  wire   [7:0] top_AND_M54_U1_t_reg;
  wire   [7:0] top_AND_M54_U1_t;
  wire   [7:0] top_AND_M54_U1_OperationInst_q;
  wire   [7:0] top_AND_M55_U1_t_reg;
  wire   [7:0] top_AND_M55_U1_t;
  wire   [7:0] top_AND_M55_U1_OperationInst_q;
  wire   [7:0] top_AND_M56_U1_t_reg;
  wire   [7:0] top_AND_M56_U1_t;
  wire   [7:0] top_AND_M56_U1_OperationInst_q;
  wire   [7:0] top_AND_M57_U1_t_reg;
  wire   [7:0] top_AND_M57_U1_t;
  wire   [7:0] top_AND_M57_U1_OperationInst_q;
  wire   [7:0] top_AND_M58_U1_t_reg;
  wire   [7:0] top_AND_M58_U1_t;
  wire   [7:0] top_AND_M58_U1_OperationInst_q;
  wire   [7:0] top_AND_M59_U1_t_reg;
  wire   [7:0] top_AND_M59_U1_t;
  wire   [7:0] top_AND_M59_U1_OperationInst_q;
  wire   [7:0] top_AND_M60_U1_t_reg;
  wire   [7:0] top_AND_M60_U1_t;
  wire   [7:0] top_AND_M60_U1_OperationInst_q;
  wire   [7:0] top_AND_M61_U1_t_reg;
  wire   [7:0] top_AND_M61_U1_t;
  wire   [7:0] top_AND_M61_U1_OperationInst_q;
  wire   [7:0] top_AND_M62_U1_t_reg;
  wire   [7:0] top_AND_M62_U1_t;
  wire   [7:0] top_AND_M62_U1_OperationInst_q;
  wire   [7:0] top_AND_M63_U1_t_reg;
  wire   [7:0] top_AND_M63_U1_t;
  wire   [7:0] top_AND_M63_U1_OperationInst_q;
  wire   [3:0] top_XOR_L0_U1_w;
  wire   [3:0] top_XOR_L1_U1_w;
  wire   [3:0] top_XOR_L2_U1_w;
  wire   [3:0] top_XOR_L3_U1_w;
  wire   [3:0] top_XOR_L4_U1_w;
  wire   [3:0] top_XOR_L5_U1_w;
  wire   [3:0] top_XOR_L6_U1_w;
  wire   [3:0] top_XOR_L7_U1_w;
  wire   [3:0] top_XOR_L8_U1_w;
  wire   [3:0] top_XOR_L9_U1_w;
  wire   [3:0] top_XOR_L10_U1_w;
  wire   [3:0] top_XOR_L11_U1_w;
  wire   [3:0] top_XOR_L12_U1_w;
  wire   [3:0] top_XOR_L13_U1_w;
  wire   [3:0] top_XOR_L14_U1_w;
  wire   [3:0] top_XOR_L15_U1_w;
  wire   [3:0] top_XOR_L16_U1_w;
  wire   [3:0] top_XOR_L17_U1_w;
  wire   [3:0] top_XOR_L18_U1_w;
  wire   [3:0] top_XOR_L19_U1_w;
  wire   [3:0] top_XOR_L20_U1_w;
  wire   [3:0] top_XOR_L21_U1_w;
  wire   [3:0] top_XOR_L22_U1_w;
  wire   [3:0] top_XOR_L23_U1_w;
  wire   [3:0] top_XOR_L24_U1_w;
  wire   [3:0] top_XOR_L25_U1_w;
  wire   [3:0] top_XOR_L26_U1_w;
  wire   [3:0] top_XOR_L27_U1_w;
  wire   [3:0] top_XOR_L28_U1_w;
  wire   [3:0] top_XOR_L29_U1_w;
  wire   [3:0] top_XOR_S0_U1_w;
  wire   [3:0] top_XOR_S1_U1_w;
  wire   [3:0] top_XOR_S2_U1_w;
  wire   [3:0] top_XOR_S3_U1_w;
  wire   [3:0] top_XOR_S4_U1_w;
  wire   [3:0] top_XOR_S5_U1_w;
  wire   [3:0] top_XOR_S6_U1_w;
  wire   [3:0] top_XOR_S7_U1_w;

  INV_X1 top_XOR_T1_U1_xorInst_U5 ( .A(top_XOR_T1_U1_xorInst_n2), .ZN(
        top_XOR_T1_U1_xorInst_n3) );
  OR2_X1 top_XOR_T1_U1_xorInst_U4 ( .A1(top_XOR_T1_U1_xorInst_n1), .A2(X_s0[7]), .ZN(top_XOR_T1_U1_xorInst_n2) );
  AND2_X1 top_XOR_T1_U1_xorInst_U3 ( .A1(X_s0[7]), .A2(
        top_XOR_T1_U1_xorInst_n1), .ZN(top_XOR_T1_U1_xorInst_n4) );
  INV_X1 top_XOR_T1_U1_xorInst_U2 ( .A(X_s0[4]), .ZN(top_XOR_T1_U1_xorInst_n1)
         );
  OR2_X1 top_XOR_T1_U1_xorInst_U1 ( .A1(top_XOR_T1_U1_xorInst_n4), .A2(
        top_XOR_T1_U1_xorInst_n3), .ZN(top_T1) );
  AND2_X1 top_XOR_T1_U1_andInst0_U1 ( .A1(X_s1[4]), .A2(X_s1_bar[7]), .ZN(
        top_XOR_T1_U1_w[0]) );
  AND2_X1 top_XOR_T1_U1_andInst1_U1 ( .A1(X_s1_bar[4]), .A2(X_s1[7]), .ZN(
        top_XOR_T1_U1_w[1]) );
  AND2_X1 top_XOR_T1_U1_andInst2_U1 ( .A1(X_s1_bar[4]), .A2(X_s1_bar[7]), .ZN(
        top_XOR_T1_U1_w[2]) );
  AND2_X1 top_XOR_T1_U1_andInst3_U1 ( .A1(X_s1[4]), .A2(X_s1[7]), .ZN(
        top_XOR_T1_U1_w[3]) );
  OR2_X1 top_XOR_T1_U1_orInst1_U1 ( .A1(top_XOR_T1_U1_w[0]), .A2(
        top_XOR_T1_U1_w[1]), .ZN(top_new_AGEMA_signal_159) );
  OR2_X1 top_XOR_T1_U1_orInst2_U1 ( .A1(top_XOR_T1_U1_w[2]), .A2(
        top_XOR_T1_U1_w[3]), .ZN(top_new_AGEMA_signal_160) );
  OR2_X1 top_XOR_T2_U1_xorInst_U5 ( .A1(top_XOR_T2_U1_xorInst_n12), .A2(
        top_XOR_T2_U1_xorInst_n11), .ZN(top_T2) );
  INV_X1 top_XOR_T2_U1_xorInst_U4 ( .A(top_XOR_T2_U1_xorInst_n10), .ZN(
        top_XOR_T2_U1_xorInst_n11) );
  OR2_X1 top_XOR_T2_U1_xorInst_U3 ( .A1(top_XOR_T2_U1_xorInst_n9), .A2(X_s0[7]), .ZN(top_XOR_T2_U1_xorInst_n10) );
  AND2_X1 top_XOR_T2_U1_xorInst_U2 ( .A1(X_s0[7]), .A2(
        top_XOR_T2_U1_xorInst_n9), .ZN(top_XOR_T2_U1_xorInst_n12) );
  INV_X1 top_XOR_T2_U1_xorInst_U1 ( .A(X_s0[2]), .ZN(top_XOR_T2_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_T2_U1_andInst0_U1 ( .A1(X_s1[2]), .A2(X_s1_bar[7]), .ZN(
        top_XOR_T2_U1_w[0]) );
  AND2_X1 top_XOR_T2_U1_andInst1_U1 ( .A1(X_s1_bar[2]), .A2(X_s1[7]), .ZN(
        top_XOR_T2_U1_w[1]) );
  AND2_X1 top_XOR_T2_U1_andInst2_U1 ( .A1(X_s1_bar[2]), .A2(X_s1_bar[7]), .ZN(
        top_XOR_T2_U1_w[2]) );
  AND2_X1 top_XOR_T2_U1_andInst3_U1 ( .A1(X_s1[2]), .A2(X_s1[7]), .ZN(
        top_XOR_T2_U1_w[3]) );
  OR2_X1 top_XOR_T2_U1_orInst1_U1 ( .A1(top_XOR_T2_U1_w[0]), .A2(
        top_XOR_T2_U1_w[1]), .ZN(top_new_AGEMA_signal_163) );
  OR2_X1 top_XOR_T2_U1_orInst2_U1 ( .A1(top_XOR_T2_U1_w[2]), .A2(
        top_XOR_T2_U1_w[3]), .ZN(top_new_AGEMA_signal_164) );
  OR2_X1 top_XOR_T3_U1_xorInst_U5 ( .A1(top_XOR_T3_U1_xorInst_n12), .A2(
        top_XOR_T3_U1_xorInst_n11), .ZN(top_T3) );
  INV_X1 top_XOR_T3_U1_xorInst_U4 ( .A(top_XOR_T3_U1_xorInst_n10), .ZN(
        top_XOR_T3_U1_xorInst_n11) );
  OR2_X1 top_XOR_T3_U1_xorInst_U3 ( .A1(top_XOR_T3_U1_xorInst_n9), .A2(X_s0[7]), .ZN(top_XOR_T3_U1_xorInst_n10) );
  AND2_X1 top_XOR_T3_U1_xorInst_U2 ( .A1(X_s0[7]), .A2(
        top_XOR_T3_U1_xorInst_n9), .ZN(top_XOR_T3_U1_xorInst_n12) );
  INV_X1 top_XOR_T3_U1_xorInst_U1 ( .A(X_s0[1]), .ZN(top_XOR_T3_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_T3_U1_andInst0_U1 ( .A1(X_s1[1]), .A2(X_s1_bar[7]), .ZN(
        top_XOR_T3_U1_w[0]) );
  AND2_X1 top_XOR_T3_U1_andInst1_U1 ( .A1(X_s1_bar[1]), .A2(X_s1[7]), .ZN(
        top_XOR_T3_U1_w[1]) );
  AND2_X1 top_XOR_T3_U1_andInst2_U1 ( .A1(X_s1_bar[1]), .A2(X_s1_bar[7]), .ZN(
        top_XOR_T3_U1_w[2]) );
  AND2_X1 top_XOR_T3_U1_andInst3_U1 ( .A1(X_s1[1]), .A2(X_s1[7]), .ZN(
        top_XOR_T3_U1_w[3]) );
  OR2_X1 top_XOR_T3_U1_orInst1_U1 ( .A1(top_XOR_T3_U1_w[0]), .A2(
        top_XOR_T3_U1_w[1]), .ZN(top_new_AGEMA_signal_167) );
  OR2_X1 top_XOR_T3_U1_orInst2_U1 ( .A1(top_XOR_T3_U1_w[2]), .A2(
        top_XOR_T3_U1_w[3]), .ZN(top_new_AGEMA_signal_168) );
  OR2_X1 top_XOR_T4_U1_xorInst_U5 ( .A1(top_XOR_T4_U1_xorInst_n12), .A2(
        top_XOR_T4_U1_xorInst_n11), .ZN(top_T4) );
  INV_X1 top_XOR_T4_U1_xorInst_U4 ( .A(top_XOR_T4_U1_xorInst_n10), .ZN(
        top_XOR_T4_U1_xorInst_n11) );
  OR2_X1 top_XOR_T4_U1_xorInst_U3 ( .A1(top_XOR_T4_U1_xorInst_n9), .A2(X_s0[4]), .ZN(top_XOR_T4_U1_xorInst_n10) );
  AND2_X1 top_XOR_T4_U1_xorInst_U2 ( .A1(X_s0[4]), .A2(
        top_XOR_T4_U1_xorInst_n9), .ZN(top_XOR_T4_U1_xorInst_n12) );
  INV_X1 top_XOR_T4_U1_xorInst_U1 ( .A(X_s0[2]), .ZN(top_XOR_T4_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_T4_U1_andInst0_U1 ( .A1(X_s1[2]), .A2(X_s1_bar[4]), .ZN(
        top_XOR_T4_U1_w[0]) );
  AND2_X1 top_XOR_T4_U1_andInst1_U1 ( .A1(X_s1_bar[2]), .A2(X_s1[4]), .ZN(
        top_XOR_T4_U1_w[1]) );
  AND2_X1 top_XOR_T4_U1_andInst2_U1 ( .A1(X_s1_bar[2]), .A2(X_s1_bar[4]), .ZN(
        top_XOR_T4_U1_w[2]) );
  AND2_X1 top_XOR_T4_U1_andInst3_U1 ( .A1(X_s1[2]), .A2(X_s1[4]), .ZN(
        top_XOR_T4_U1_w[3]) );
  OR2_X1 top_XOR_T4_U1_orInst1_U1 ( .A1(top_XOR_T4_U1_w[0]), .A2(
        top_XOR_T4_U1_w[1]), .ZN(top_new_AGEMA_signal_169) );
  OR2_X1 top_XOR_T4_U1_orInst2_U1 ( .A1(top_XOR_T4_U1_w[2]), .A2(
        top_XOR_T4_U1_w[3]), .ZN(top_new_AGEMA_signal_170) );
  OR2_X1 top_XOR_T5_U1_xorInst_U5 ( .A1(top_XOR_T5_U1_xorInst_n12), .A2(
        top_XOR_T5_U1_xorInst_n11), .ZN(top_T5) );
  INV_X1 top_XOR_T5_U1_xorInst_U4 ( .A(top_XOR_T5_U1_xorInst_n10), .ZN(
        top_XOR_T5_U1_xorInst_n11) );
  OR2_X1 top_XOR_T5_U1_xorInst_U3 ( .A1(top_XOR_T5_U1_xorInst_n9), .A2(X_s0[3]), .ZN(top_XOR_T5_U1_xorInst_n10) );
  AND2_X1 top_XOR_T5_U1_xorInst_U2 ( .A1(X_s0[3]), .A2(
        top_XOR_T5_U1_xorInst_n9), .ZN(top_XOR_T5_U1_xorInst_n12) );
  INV_X1 top_XOR_T5_U1_xorInst_U1 ( .A(X_s0[1]), .ZN(top_XOR_T5_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_T5_U1_andInst0_U1 ( .A1(X_s1[1]), .A2(X_s1_bar[3]), .ZN(
        top_XOR_T5_U1_w[0]) );
  AND2_X1 top_XOR_T5_U1_andInst1_U1 ( .A1(X_s1_bar[1]), .A2(X_s1[3]), .ZN(
        top_XOR_T5_U1_w[1]) );
  AND2_X1 top_XOR_T5_U1_andInst2_U1 ( .A1(X_s1_bar[1]), .A2(X_s1_bar[3]), .ZN(
        top_XOR_T5_U1_w[2]) );
  AND2_X1 top_XOR_T5_U1_andInst3_U1 ( .A1(X_s1[1]), .A2(X_s1[3]), .ZN(
        top_XOR_T5_U1_w[3]) );
  OR2_X1 top_XOR_T5_U1_orInst1_U1 ( .A1(top_XOR_T5_U1_w[0]), .A2(
        top_XOR_T5_U1_w[1]), .ZN(top_new_AGEMA_signal_173) );
  OR2_X1 top_XOR_T5_U1_orInst2_U1 ( .A1(top_XOR_T5_U1_w[2]), .A2(
        top_XOR_T5_U1_w[3]), .ZN(top_new_AGEMA_signal_174) );
  OR2_X1 top_XOR_T6_U1_xorInst_U5 ( .A1(top_XOR_T6_U1_xorInst_n12), .A2(
        top_XOR_T6_U1_xorInst_n11), .ZN(top_T6) );
  INV_X1 top_XOR_T6_U1_xorInst_U4 ( .A(top_XOR_T6_U1_xorInst_n10), .ZN(
        top_XOR_T6_U1_xorInst_n11) );
  OR2_X1 top_XOR_T6_U1_xorInst_U3 ( .A1(top_XOR_T6_U1_xorInst_n9), .A2(top_T1), 
        .ZN(top_XOR_T6_U1_xorInst_n10) );
  AND2_X1 top_XOR_T6_U1_xorInst_U2 ( .A1(top_T1), .A2(top_XOR_T6_U1_xorInst_n9), .ZN(top_XOR_T6_U1_xorInst_n12) );
  INV_X1 top_XOR_T6_U1_xorInst_U1 ( .A(top_T5), .ZN(top_XOR_T6_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_T6_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_173), .A2(
        top_new_AGEMA_signal_160), .ZN(top_XOR_T6_U1_w[0]) );
  AND2_X1 top_XOR_T6_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_174), .A2(
        top_new_AGEMA_signal_159), .ZN(top_XOR_T6_U1_w[1]) );
  AND2_X1 top_XOR_T6_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_174), .A2(
        top_new_AGEMA_signal_160), .ZN(top_XOR_T6_U1_w[2]) );
  AND2_X1 top_XOR_T6_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_173), .A2(
        top_new_AGEMA_signal_159), .ZN(top_XOR_T6_U1_w[3]) );
  OR2_X1 top_XOR_T6_U1_orInst1_U1 ( .A1(top_XOR_T6_U1_w[0]), .A2(
        top_XOR_T6_U1_w[1]), .ZN(top_new_AGEMA_signal_191) );
  OR2_X1 top_XOR_T6_U1_orInst2_U1 ( .A1(top_XOR_T6_U1_w[2]), .A2(
        top_XOR_T6_U1_w[3]), .ZN(top_new_AGEMA_signal_192) );
  OR2_X1 top_XOR_T7_U1_xorInst_U5 ( .A1(top_XOR_T7_U1_xorInst_n12), .A2(
        top_XOR_T7_U1_xorInst_n11), .ZN(top_T7) );
  INV_X1 top_XOR_T7_U1_xorInst_U4 ( .A(top_XOR_T7_U1_xorInst_n10), .ZN(
        top_XOR_T7_U1_xorInst_n11) );
  OR2_X1 top_XOR_T7_U1_xorInst_U3 ( .A1(top_XOR_T7_U1_xorInst_n9), .A2(X_s0[6]), .ZN(top_XOR_T7_U1_xorInst_n10) );
  AND2_X1 top_XOR_T7_U1_xorInst_U2 ( .A1(X_s0[6]), .A2(
        top_XOR_T7_U1_xorInst_n9), .ZN(top_XOR_T7_U1_xorInst_n12) );
  INV_X1 top_XOR_T7_U1_xorInst_U1 ( .A(X_s0[5]), .ZN(top_XOR_T7_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_T7_U1_andInst0_U1 ( .A1(X_s1[5]), .A2(X_s1_bar[6]), .ZN(
        top_XOR_T7_U1_w[0]) );
  AND2_X1 top_XOR_T7_U1_andInst1_U1 ( .A1(X_s1_bar[5]), .A2(X_s1[6]), .ZN(
        top_XOR_T7_U1_w[1]) );
  AND2_X1 top_XOR_T7_U1_andInst2_U1 ( .A1(X_s1_bar[5]), .A2(X_s1_bar[6]), .ZN(
        top_XOR_T7_U1_w[2]) );
  AND2_X1 top_XOR_T7_U1_andInst3_U1 ( .A1(X_s1[5]), .A2(X_s1[6]), .ZN(
        top_XOR_T7_U1_w[3]) );
  OR2_X1 top_XOR_T7_U1_orInst1_U1 ( .A1(top_XOR_T7_U1_w[0]), .A2(
        top_XOR_T7_U1_w[1]), .ZN(top_new_AGEMA_signal_179) );
  OR2_X1 top_XOR_T7_U1_orInst2_U1 ( .A1(top_XOR_T7_U1_w[2]), .A2(
        top_XOR_T7_U1_w[3]), .ZN(top_new_AGEMA_signal_180) );
  OR2_X1 top_XOR_T8_U1_xorInst_U5 ( .A1(top_XOR_T8_U1_xorInst_n12), .A2(
        top_XOR_T8_U1_xorInst_n11), .ZN(top_T8) );
  INV_X1 top_XOR_T8_U1_xorInst_U4 ( .A(top_XOR_T8_U1_xorInst_n10), .ZN(
        top_XOR_T8_U1_xorInst_n11) );
  OR2_X1 top_XOR_T8_U1_xorInst_U3 ( .A1(top_XOR_T8_U1_xorInst_n9), .A2(X_s0[0]), .ZN(top_XOR_T8_U1_xorInst_n10) );
  AND2_X1 top_XOR_T8_U1_xorInst_U2 ( .A1(X_s0[0]), .A2(
        top_XOR_T8_U1_xorInst_n9), .ZN(top_XOR_T8_U1_xorInst_n12) );
  INV_X1 top_XOR_T8_U1_xorInst_U1 ( .A(top_T6), .ZN(top_XOR_T8_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_T8_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_191), .A2(
        X_s1_bar[0]), .ZN(top_XOR_T8_U1_w[0]) );
  AND2_X1 top_XOR_T8_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_192), .A2(
        X_s1[0]), .ZN(top_XOR_T8_U1_w[1]) );
  AND2_X1 top_XOR_T8_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_192), .A2(
        X_s1_bar[0]), .ZN(top_XOR_T8_U1_w[2]) );
  AND2_X1 top_XOR_T8_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_191), .A2(
        X_s1[0]), .ZN(top_XOR_T8_U1_w[3]) );
  OR2_X1 top_XOR_T8_U1_orInst1_U1 ( .A1(top_XOR_T8_U1_w[0]), .A2(
        top_XOR_T8_U1_w[1]), .ZN(top_new_AGEMA_signal_207) );
  OR2_X1 top_XOR_T8_U1_orInst2_U1 ( .A1(top_XOR_T8_U1_w[2]), .A2(
        top_XOR_T8_U1_w[3]), .ZN(top_new_AGEMA_signal_208) );
  OR2_X1 top_XOR_T9_U1_xorInst_U5 ( .A1(top_XOR_T9_U1_xorInst_n12), .A2(
        top_XOR_T9_U1_xorInst_n11), .ZN(top_T9) );
  INV_X1 top_XOR_T9_U1_xorInst_U4 ( .A(top_XOR_T9_U1_xorInst_n10), .ZN(
        top_XOR_T9_U1_xorInst_n11) );
  OR2_X1 top_XOR_T9_U1_xorInst_U3 ( .A1(top_XOR_T9_U1_xorInst_n9), .A2(X_s0[0]), .ZN(top_XOR_T9_U1_xorInst_n10) );
  AND2_X1 top_XOR_T9_U1_xorInst_U2 ( .A1(X_s0[0]), .A2(
        top_XOR_T9_U1_xorInst_n9), .ZN(top_XOR_T9_U1_xorInst_n12) );
  INV_X1 top_XOR_T9_U1_xorInst_U1 ( .A(top_T7), .ZN(top_XOR_T9_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_T9_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_179), .A2(
        X_s1_bar[0]), .ZN(top_XOR_T9_U1_w[0]) );
  AND2_X1 top_XOR_T9_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_180), .A2(
        X_s1[0]), .ZN(top_XOR_T9_U1_w[1]) );
  AND2_X1 top_XOR_T9_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_180), .A2(
        X_s1_bar[0]), .ZN(top_XOR_T9_U1_w[2]) );
  AND2_X1 top_XOR_T9_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_179), .A2(
        X_s1[0]), .ZN(top_XOR_T9_U1_w[3]) );
  OR2_X1 top_XOR_T9_U1_orInst1_U1 ( .A1(top_XOR_T9_U1_w[0]), .A2(
        top_XOR_T9_U1_w[1]), .ZN(top_new_AGEMA_signal_193) );
  OR2_X1 top_XOR_T9_U1_orInst2_U1 ( .A1(top_XOR_T9_U1_w[2]), .A2(
        top_XOR_T9_U1_w[3]), .ZN(top_new_AGEMA_signal_194) );
  OR2_X1 top_XOR_T10_U1_xorInst_U5 ( .A1(top_XOR_T10_U1_xorInst_n12), .A2(
        top_XOR_T10_U1_xorInst_n11), .ZN(top_T10) );
  INV_X1 top_XOR_T10_U1_xorInst_U4 ( .A(top_XOR_T10_U1_xorInst_n10), .ZN(
        top_XOR_T10_U1_xorInst_n11) );
  OR2_X1 top_XOR_T10_U1_xorInst_U3 ( .A1(top_XOR_T10_U1_xorInst_n9), .A2(
        top_T6), .ZN(top_XOR_T10_U1_xorInst_n10) );
  AND2_X1 top_XOR_T10_U1_xorInst_U2 ( .A1(top_T6), .A2(
        top_XOR_T10_U1_xorInst_n9), .ZN(top_XOR_T10_U1_xorInst_n12) );
  INV_X1 top_XOR_T10_U1_xorInst_U1 ( .A(top_T7), .ZN(top_XOR_T10_U1_xorInst_n9) );
  AND2_X1 top_XOR_T10_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_179), .A2(
        top_new_AGEMA_signal_192), .ZN(top_XOR_T10_U1_w[0]) );
  AND2_X1 top_XOR_T10_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_180), .A2(
        top_new_AGEMA_signal_191), .ZN(top_XOR_T10_U1_w[1]) );
  AND2_X1 top_XOR_T10_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_180), .A2(
        top_new_AGEMA_signal_192), .ZN(top_XOR_T10_U1_w[2]) );
  AND2_X1 top_XOR_T10_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_179), .A2(
        top_new_AGEMA_signal_191), .ZN(top_XOR_T10_U1_w[3]) );
  OR2_X1 top_XOR_T10_U1_orInst1_U1 ( .A1(top_XOR_T10_U1_w[0]), .A2(
        top_XOR_T10_U1_w[1]), .ZN(top_new_AGEMA_signal_209) );
  OR2_X1 top_XOR_T10_U1_orInst2_U1 ( .A1(top_XOR_T10_U1_w[2]), .A2(
        top_XOR_T10_U1_w[3]), .ZN(top_new_AGEMA_signal_210) );
  OR2_X1 top_XOR_T11_U1_xorInst_U5 ( .A1(top_XOR_T11_U1_xorInst_n12), .A2(
        top_XOR_T11_U1_xorInst_n11), .ZN(top_T11) );
  INV_X1 top_XOR_T11_U1_xorInst_U4 ( .A(top_XOR_T11_U1_xorInst_n10), .ZN(
        top_XOR_T11_U1_xorInst_n11) );
  OR2_X1 top_XOR_T11_U1_xorInst_U3 ( .A1(top_XOR_T11_U1_xorInst_n9), .A2(
        X_s0[6]), .ZN(top_XOR_T11_U1_xorInst_n10) );
  AND2_X1 top_XOR_T11_U1_xorInst_U2 ( .A1(X_s0[6]), .A2(
        top_XOR_T11_U1_xorInst_n9), .ZN(top_XOR_T11_U1_xorInst_n12) );
  INV_X1 top_XOR_T11_U1_xorInst_U1 ( .A(X_s0[2]), .ZN(
        top_XOR_T11_U1_xorInst_n9) );
  AND2_X1 top_XOR_T11_U1_andInst0_U1 ( .A1(X_s1[2]), .A2(X_s1_bar[6]), .ZN(
        top_XOR_T11_U1_w[0]) );
  AND2_X1 top_XOR_T11_U1_andInst1_U1 ( .A1(X_s1_bar[2]), .A2(X_s1[6]), .ZN(
        top_XOR_T11_U1_w[1]) );
  AND2_X1 top_XOR_T11_U1_andInst2_U1 ( .A1(X_s1_bar[2]), .A2(X_s1_bar[6]), 
        .ZN(top_XOR_T11_U1_w[2]) );
  AND2_X1 top_XOR_T11_U1_andInst3_U1 ( .A1(X_s1[2]), .A2(X_s1[6]), .ZN(
        top_XOR_T11_U1_w[3]) );
  OR2_X1 top_XOR_T11_U1_orInst1_U1 ( .A1(top_XOR_T11_U1_w[0]), .A2(
        top_XOR_T11_U1_w[1]), .ZN(top_new_AGEMA_signal_181) );
  OR2_X1 top_XOR_T11_U1_orInst2_U1 ( .A1(top_XOR_T11_U1_w[2]), .A2(
        top_XOR_T11_U1_w[3]), .ZN(top_new_AGEMA_signal_182) );
  OR2_X1 top_XOR_T12_U1_xorInst_U5 ( .A1(top_XOR_T12_U1_xorInst_n12), .A2(
        top_XOR_T12_U1_xorInst_n11), .ZN(top_T12) );
  INV_X1 top_XOR_T12_U1_xorInst_U4 ( .A(top_XOR_T12_U1_xorInst_n10), .ZN(
        top_XOR_T12_U1_xorInst_n11) );
  OR2_X1 top_XOR_T12_U1_xorInst_U3 ( .A1(top_XOR_T12_U1_xorInst_n9), .A2(
        X_s0[5]), .ZN(top_XOR_T12_U1_xorInst_n10) );
  AND2_X1 top_XOR_T12_U1_xorInst_U2 ( .A1(X_s0[5]), .A2(
        top_XOR_T12_U1_xorInst_n9), .ZN(top_XOR_T12_U1_xorInst_n12) );
  INV_X1 top_XOR_T12_U1_xorInst_U1 ( .A(X_s0[2]), .ZN(
        top_XOR_T12_U1_xorInst_n9) );
  AND2_X1 top_XOR_T12_U1_andInst0_U1 ( .A1(X_s1[2]), .A2(X_s1_bar[5]), .ZN(
        top_XOR_T12_U1_w[0]) );
  AND2_X1 top_XOR_T12_U1_andInst1_U1 ( .A1(X_s1_bar[2]), .A2(X_s1[5]), .ZN(
        top_XOR_T12_U1_w[1]) );
  AND2_X1 top_XOR_T12_U1_andInst2_U1 ( .A1(X_s1_bar[2]), .A2(X_s1_bar[5]), 
        .ZN(top_XOR_T12_U1_w[2]) );
  AND2_X1 top_XOR_T12_U1_andInst3_U1 ( .A1(X_s1[2]), .A2(X_s1[5]), .ZN(
        top_XOR_T12_U1_w[3]) );
  OR2_X1 top_XOR_T12_U1_orInst1_U1 ( .A1(top_XOR_T12_U1_w[0]), .A2(
        top_XOR_T12_U1_w[1]), .ZN(top_new_AGEMA_signal_183) );
  OR2_X1 top_XOR_T12_U1_orInst2_U1 ( .A1(top_XOR_T12_U1_w[2]), .A2(
        top_XOR_T12_U1_w[3]), .ZN(top_new_AGEMA_signal_184) );
  OR2_X1 top_XOR_T13_U1_xorInst_U5 ( .A1(top_XOR_T13_U1_xorInst_n12), .A2(
        top_XOR_T13_U1_xorInst_n11), .ZN(top_T13) );
  INV_X1 top_XOR_T13_U1_xorInst_U4 ( .A(top_XOR_T13_U1_xorInst_n10), .ZN(
        top_XOR_T13_U1_xorInst_n11) );
  OR2_X1 top_XOR_T13_U1_xorInst_U3 ( .A1(top_XOR_T13_U1_xorInst_n9), .A2(
        top_T3), .ZN(top_XOR_T13_U1_xorInst_n10) );
  AND2_X1 top_XOR_T13_U1_xorInst_U2 ( .A1(top_T3), .A2(
        top_XOR_T13_U1_xorInst_n9), .ZN(top_XOR_T13_U1_xorInst_n12) );
  INV_X1 top_XOR_T13_U1_xorInst_U1 ( .A(top_T4), .ZN(top_XOR_T13_U1_xorInst_n9) );
  AND2_X1 top_XOR_T13_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_169), .A2(
        top_new_AGEMA_signal_168), .ZN(top_XOR_T13_U1_w[0]) );
  AND2_X1 top_XOR_T13_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_170), .A2(
        top_new_AGEMA_signal_167), .ZN(top_XOR_T13_U1_w[1]) );
  AND2_X1 top_XOR_T13_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_170), .A2(
        top_new_AGEMA_signal_168), .ZN(top_XOR_T13_U1_w[2]) );
  AND2_X1 top_XOR_T13_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_169), .A2(
        top_new_AGEMA_signal_167), .ZN(top_XOR_T13_U1_w[3]) );
  OR2_X1 top_XOR_T13_U1_orInst1_U1 ( .A1(top_XOR_T13_U1_w[0]), .A2(
        top_XOR_T13_U1_w[1]), .ZN(top_new_AGEMA_signal_195) );
  OR2_X1 top_XOR_T13_U1_orInst2_U1 ( .A1(top_XOR_T13_U1_w[2]), .A2(
        top_XOR_T13_U1_w[3]), .ZN(top_new_AGEMA_signal_196) );
  OR2_X1 top_XOR_T14_U1_xorInst_U5 ( .A1(top_XOR_T14_U1_xorInst_n12), .A2(
        top_XOR_T14_U1_xorInst_n11), .ZN(top_T14) );
  INV_X1 top_XOR_T14_U1_xorInst_U4 ( .A(top_XOR_T14_U1_xorInst_n10), .ZN(
        top_XOR_T14_U1_xorInst_n11) );
  OR2_X1 top_XOR_T14_U1_xorInst_U3 ( .A1(top_XOR_T14_U1_xorInst_n9), .A2(
        top_T6), .ZN(top_XOR_T14_U1_xorInst_n10) );
  AND2_X1 top_XOR_T14_U1_xorInst_U2 ( .A1(top_T6), .A2(
        top_XOR_T14_U1_xorInst_n9), .ZN(top_XOR_T14_U1_xorInst_n12) );
  INV_X1 top_XOR_T14_U1_xorInst_U1 ( .A(top_T11), .ZN(
        top_XOR_T14_U1_xorInst_n9) );
  AND2_X1 top_XOR_T14_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_181), .A2(
        top_new_AGEMA_signal_192), .ZN(top_XOR_T14_U1_w[0]) );
  AND2_X1 top_XOR_T14_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_182), .A2(
        top_new_AGEMA_signal_191), .ZN(top_XOR_T14_U1_w[1]) );
  AND2_X1 top_XOR_T14_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_182), .A2(
        top_new_AGEMA_signal_192), .ZN(top_XOR_T14_U1_w[2]) );
  AND2_X1 top_XOR_T14_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_181), .A2(
        top_new_AGEMA_signal_191), .ZN(top_XOR_T14_U1_w[3]) );
  OR2_X1 top_XOR_T14_U1_orInst1_U1 ( .A1(top_XOR_T14_U1_w[0]), .A2(
        top_XOR_T14_U1_w[1]), .ZN(top_new_AGEMA_signal_211) );
  OR2_X1 top_XOR_T14_U1_orInst2_U1 ( .A1(top_XOR_T14_U1_w[2]), .A2(
        top_XOR_T14_U1_w[3]), .ZN(top_new_AGEMA_signal_212) );
  OR2_X1 top_XOR_T15_U1_xorInst_U5 ( .A1(top_XOR_T15_U1_xorInst_n12), .A2(
        top_XOR_T15_U1_xorInst_n11), .ZN(top_T15) );
  INV_X1 top_XOR_T15_U1_xorInst_U4 ( .A(top_XOR_T15_U1_xorInst_n10), .ZN(
        top_XOR_T15_U1_xorInst_n11) );
  OR2_X1 top_XOR_T15_U1_xorInst_U3 ( .A1(top_XOR_T15_U1_xorInst_n9), .A2(
        top_T5), .ZN(top_XOR_T15_U1_xorInst_n10) );
  AND2_X1 top_XOR_T15_U1_xorInst_U2 ( .A1(top_T5), .A2(
        top_XOR_T15_U1_xorInst_n9), .ZN(top_XOR_T15_U1_xorInst_n12) );
  INV_X1 top_XOR_T15_U1_xorInst_U1 ( .A(top_T11), .ZN(
        top_XOR_T15_U1_xorInst_n9) );
  AND2_X1 top_XOR_T15_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_181), .A2(
        top_new_AGEMA_signal_174), .ZN(top_XOR_T15_U1_w[0]) );
  AND2_X1 top_XOR_T15_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_182), .A2(
        top_new_AGEMA_signal_173), .ZN(top_XOR_T15_U1_w[1]) );
  AND2_X1 top_XOR_T15_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_182), .A2(
        top_new_AGEMA_signal_174), .ZN(top_XOR_T15_U1_w[2]) );
  AND2_X1 top_XOR_T15_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_181), .A2(
        top_new_AGEMA_signal_173), .ZN(top_XOR_T15_U1_w[3]) );
  OR2_X1 top_XOR_T15_U1_orInst1_U1 ( .A1(top_XOR_T15_U1_w[0]), .A2(
        top_XOR_T15_U1_w[1]), .ZN(top_new_AGEMA_signal_197) );
  OR2_X1 top_XOR_T15_U1_orInst2_U1 ( .A1(top_XOR_T15_U1_w[2]), .A2(
        top_XOR_T15_U1_w[3]), .ZN(top_new_AGEMA_signal_198) );
  OR2_X1 top_XOR_T16_U1_xorInst_U5 ( .A1(top_XOR_T16_U1_xorInst_n12), .A2(
        top_XOR_T16_U1_xorInst_n11), .ZN(top_T16) );
  INV_X1 top_XOR_T16_U1_xorInst_U4 ( .A(top_XOR_T16_U1_xorInst_n10), .ZN(
        top_XOR_T16_U1_xorInst_n11) );
  OR2_X1 top_XOR_T16_U1_xorInst_U3 ( .A1(top_XOR_T16_U1_xorInst_n9), .A2(
        top_T5), .ZN(top_XOR_T16_U1_xorInst_n10) );
  AND2_X1 top_XOR_T16_U1_xorInst_U2 ( .A1(top_T5), .A2(
        top_XOR_T16_U1_xorInst_n9), .ZN(top_XOR_T16_U1_xorInst_n12) );
  INV_X1 top_XOR_T16_U1_xorInst_U1 ( .A(top_T12), .ZN(
        top_XOR_T16_U1_xorInst_n9) );
  AND2_X1 top_XOR_T16_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_183), .A2(
        top_new_AGEMA_signal_174), .ZN(top_XOR_T16_U1_w[0]) );
  AND2_X1 top_XOR_T16_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_184), .A2(
        top_new_AGEMA_signal_173), .ZN(top_XOR_T16_U1_w[1]) );
  AND2_X1 top_XOR_T16_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_184), .A2(
        top_new_AGEMA_signal_174), .ZN(top_XOR_T16_U1_w[2]) );
  AND2_X1 top_XOR_T16_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_183), .A2(
        top_new_AGEMA_signal_173), .ZN(top_XOR_T16_U1_w[3]) );
  OR2_X1 top_XOR_T16_U1_orInst1_U1 ( .A1(top_XOR_T16_U1_w[0]), .A2(
        top_XOR_T16_U1_w[1]), .ZN(top_new_AGEMA_signal_199) );
  OR2_X1 top_XOR_T16_U1_orInst2_U1 ( .A1(top_XOR_T16_U1_w[2]), .A2(
        top_XOR_T16_U1_w[3]), .ZN(top_new_AGEMA_signal_200) );
  OR2_X1 top_XOR_T17_U1_xorInst_U5 ( .A1(top_XOR_T17_U1_xorInst_n12), .A2(
        top_XOR_T17_U1_xorInst_n11), .ZN(top_T17) );
  INV_X1 top_XOR_T17_U1_xorInst_U4 ( .A(top_XOR_T17_U1_xorInst_n10), .ZN(
        top_XOR_T17_U1_xorInst_n11) );
  OR2_X1 top_XOR_T17_U1_xorInst_U3 ( .A1(top_XOR_T17_U1_xorInst_n9), .A2(
        top_T9), .ZN(top_XOR_T17_U1_xorInst_n10) );
  AND2_X1 top_XOR_T17_U1_xorInst_U2 ( .A1(top_T9), .A2(
        top_XOR_T17_U1_xorInst_n9), .ZN(top_XOR_T17_U1_xorInst_n12) );
  INV_X1 top_XOR_T17_U1_xorInst_U1 ( .A(top_T16), .ZN(
        top_XOR_T17_U1_xorInst_n9) );
  AND2_X1 top_XOR_T17_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_199), .A2(
        top_new_AGEMA_signal_194), .ZN(top_XOR_T17_U1_w[0]) );
  AND2_X1 top_XOR_T17_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_200), .A2(
        top_new_AGEMA_signal_193), .ZN(top_XOR_T17_U1_w[1]) );
  AND2_X1 top_XOR_T17_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_200), .A2(
        top_new_AGEMA_signal_194), .ZN(top_XOR_T17_U1_w[2]) );
  AND2_X1 top_XOR_T17_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_199), .A2(
        top_new_AGEMA_signal_193), .ZN(top_XOR_T17_U1_w[3]) );
  OR2_X1 top_XOR_T17_U1_orInst1_U1 ( .A1(top_XOR_T17_U1_w[0]), .A2(
        top_XOR_T17_U1_w[1]), .ZN(top_new_AGEMA_signal_213) );
  OR2_X1 top_XOR_T17_U1_orInst2_U1 ( .A1(top_XOR_T17_U1_w[2]), .A2(
        top_XOR_T17_U1_w[3]), .ZN(top_new_AGEMA_signal_214) );
  OR2_X1 top_XOR_T18_U1_xorInst_U5 ( .A1(top_XOR_T18_U1_xorInst_n12), .A2(
        top_XOR_T18_U1_xorInst_n11), .ZN(top_T18) );
  INV_X1 top_XOR_T18_U1_xorInst_U4 ( .A(top_XOR_T18_U1_xorInst_n10), .ZN(
        top_XOR_T18_U1_xorInst_n11) );
  OR2_X1 top_XOR_T18_U1_xorInst_U3 ( .A1(top_XOR_T18_U1_xorInst_n9), .A2(
        X_s0[4]), .ZN(top_XOR_T18_U1_xorInst_n10) );
  AND2_X1 top_XOR_T18_U1_xorInst_U2 ( .A1(X_s0[4]), .A2(
        top_XOR_T18_U1_xorInst_n9), .ZN(top_XOR_T18_U1_xorInst_n12) );
  INV_X1 top_XOR_T18_U1_xorInst_U1 ( .A(X_s0[0]), .ZN(
        top_XOR_T18_U1_xorInst_n9) );
  AND2_X1 top_XOR_T18_U1_andInst0_U1 ( .A1(X_s1[0]), .A2(X_s1_bar[4]), .ZN(
        top_XOR_T18_U1_w[0]) );
  AND2_X1 top_XOR_T18_U1_andInst1_U1 ( .A1(X_s1_bar[0]), .A2(X_s1[4]), .ZN(
        top_XOR_T18_U1_w[1]) );
  AND2_X1 top_XOR_T18_U1_andInst2_U1 ( .A1(X_s1_bar[0]), .A2(X_s1_bar[4]), 
        .ZN(top_XOR_T18_U1_w[2]) );
  AND2_X1 top_XOR_T18_U1_andInst3_U1 ( .A1(X_s1[0]), .A2(X_s1[4]), .ZN(
        top_XOR_T18_U1_w[3]) );
  OR2_X1 top_XOR_T18_U1_orInst1_U1 ( .A1(top_XOR_T18_U1_w[0]), .A2(
        top_XOR_T18_U1_w[1]), .ZN(top_new_AGEMA_signal_187) );
  OR2_X1 top_XOR_T18_U1_orInst2_U1 ( .A1(top_XOR_T18_U1_w[2]), .A2(
        top_XOR_T18_U1_w[3]), .ZN(top_new_AGEMA_signal_188) );
  OR2_X1 top_XOR_T19_U1_xorInst_U5 ( .A1(top_XOR_T19_U1_xorInst_n12), .A2(
        top_XOR_T19_U1_xorInst_n11), .ZN(top_T19) );
  INV_X1 top_XOR_T19_U1_xorInst_U4 ( .A(top_XOR_T19_U1_xorInst_n10), .ZN(
        top_XOR_T19_U1_xorInst_n11) );
  OR2_X1 top_XOR_T19_U1_xorInst_U3 ( .A1(top_XOR_T19_U1_xorInst_n9), .A2(
        top_T7), .ZN(top_XOR_T19_U1_xorInst_n10) );
  AND2_X1 top_XOR_T19_U1_xorInst_U2 ( .A1(top_T7), .A2(
        top_XOR_T19_U1_xorInst_n9), .ZN(top_XOR_T19_U1_xorInst_n12) );
  INV_X1 top_XOR_T19_U1_xorInst_U1 ( .A(top_T18), .ZN(
        top_XOR_T19_U1_xorInst_n9) );
  AND2_X1 top_XOR_T19_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_187), .A2(
        top_new_AGEMA_signal_180), .ZN(top_XOR_T19_U1_w[0]) );
  AND2_X1 top_XOR_T19_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_188), .A2(
        top_new_AGEMA_signal_179), .ZN(top_XOR_T19_U1_w[1]) );
  AND2_X1 top_XOR_T19_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_188), .A2(
        top_new_AGEMA_signal_180), .ZN(top_XOR_T19_U1_w[2]) );
  AND2_X1 top_XOR_T19_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_187), .A2(
        top_new_AGEMA_signal_179), .ZN(top_XOR_T19_U1_w[3]) );
  OR2_X1 top_XOR_T19_U1_orInst1_U1 ( .A1(top_XOR_T19_U1_w[0]), .A2(
        top_XOR_T19_U1_w[1]), .ZN(top_new_AGEMA_signal_201) );
  OR2_X1 top_XOR_T19_U1_orInst2_U1 ( .A1(top_XOR_T19_U1_w[2]), .A2(
        top_XOR_T19_U1_w[3]), .ZN(top_new_AGEMA_signal_202) );
  OR2_X1 top_XOR_T20_U1_xorInst_U5 ( .A1(top_XOR_T20_U1_xorInst_n12), .A2(
        top_XOR_T20_U1_xorInst_n11), .ZN(top_T20) );
  INV_X1 top_XOR_T20_U1_xorInst_U4 ( .A(top_XOR_T20_U1_xorInst_n10), .ZN(
        top_XOR_T20_U1_xorInst_n11) );
  OR2_X1 top_XOR_T20_U1_xorInst_U3 ( .A1(top_XOR_T20_U1_xorInst_n9), .A2(
        top_T1), .ZN(top_XOR_T20_U1_xorInst_n10) );
  AND2_X1 top_XOR_T20_U1_xorInst_U2 ( .A1(top_T1), .A2(
        top_XOR_T20_U1_xorInst_n9), .ZN(top_XOR_T20_U1_xorInst_n12) );
  INV_X1 top_XOR_T20_U1_xorInst_U1 ( .A(top_T19), .ZN(
        top_XOR_T20_U1_xorInst_n9) );
  AND2_X1 top_XOR_T20_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_201), .A2(
        top_new_AGEMA_signal_160), .ZN(top_XOR_T20_U1_w[0]) );
  AND2_X1 top_XOR_T20_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_202), .A2(
        top_new_AGEMA_signal_159), .ZN(top_XOR_T20_U1_w[1]) );
  AND2_X1 top_XOR_T20_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_202), .A2(
        top_new_AGEMA_signal_160), .ZN(top_XOR_T20_U1_w[2]) );
  AND2_X1 top_XOR_T20_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_201), .A2(
        top_new_AGEMA_signal_159), .ZN(top_XOR_T20_U1_w[3]) );
  OR2_X1 top_XOR_T20_U1_orInst1_U1 ( .A1(top_XOR_T20_U1_w[0]), .A2(
        top_XOR_T20_U1_w[1]), .ZN(top_new_AGEMA_signal_215) );
  OR2_X1 top_XOR_T20_U1_orInst2_U1 ( .A1(top_XOR_T20_U1_w[2]), .A2(
        top_XOR_T20_U1_w[3]), .ZN(top_new_AGEMA_signal_216) );
  OR2_X1 top_XOR_T21_U1_xorInst_U5 ( .A1(top_XOR_T21_U1_xorInst_n12), .A2(
        top_XOR_T21_U1_xorInst_n11), .ZN(top_T21) );
  INV_X1 top_XOR_T21_U1_xorInst_U4 ( .A(top_XOR_T21_U1_xorInst_n10), .ZN(
        top_XOR_T21_U1_xorInst_n11) );
  OR2_X1 top_XOR_T21_U1_xorInst_U3 ( .A1(top_XOR_T21_U1_xorInst_n9), .A2(
        X_s0[1]), .ZN(top_XOR_T21_U1_xorInst_n10) );
  AND2_X1 top_XOR_T21_U1_xorInst_U2 ( .A1(X_s0[1]), .A2(
        top_XOR_T21_U1_xorInst_n9), .ZN(top_XOR_T21_U1_xorInst_n12) );
  INV_X1 top_XOR_T21_U1_xorInst_U1 ( .A(X_s0[0]), .ZN(
        top_XOR_T21_U1_xorInst_n9) );
  AND2_X1 top_XOR_T21_U1_andInst0_U1 ( .A1(X_s1[0]), .A2(X_s1_bar[1]), .ZN(
        top_XOR_T21_U1_w[0]) );
  AND2_X1 top_XOR_T21_U1_andInst1_U1 ( .A1(X_s1_bar[0]), .A2(X_s1[1]), .ZN(
        top_XOR_T21_U1_w[1]) );
  AND2_X1 top_XOR_T21_U1_andInst2_U1 ( .A1(X_s1_bar[0]), .A2(X_s1_bar[1]), 
        .ZN(top_XOR_T21_U1_w[2]) );
  AND2_X1 top_XOR_T21_U1_andInst3_U1 ( .A1(X_s1[0]), .A2(X_s1[1]), .ZN(
        top_XOR_T21_U1_w[3]) );
  OR2_X1 top_XOR_T21_U1_orInst1_U1 ( .A1(top_XOR_T21_U1_w[0]), .A2(
        top_XOR_T21_U1_w[1]), .ZN(top_new_AGEMA_signal_189) );
  OR2_X1 top_XOR_T21_U1_orInst2_U1 ( .A1(top_XOR_T21_U1_w[2]), .A2(
        top_XOR_T21_U1_w[3]), .ZN(top_new_AGEMA_signal_190) );
  OR2_X1 top_XOR_T22_U1_xorInst_U5 ( .A1(top_XOR_T22_U1_xorInst_n12), .A2(
        top_XOR_T22_U1_xorInst_n11), .ZN(top_T22) );
  INV_X1 top_XOR_T22_U1_xorInst_U4 ( .A(top_XOR_T22_U1_xorInst_n10), .ZN(
        top_XOR_T22_U1_xorInst_n11) );
  OR2_X1 top_XOR_T22_U1_xorInst_U3 ( .A1(top_XOR_T22_U1_xorInst_n9), .A2(
        top_T7), .ZN(top_XOR_T22_U1_xorInst_n10) );
  AND2_X1 top_XOR_T22_U1_xorInst_U2 ( .A1(top_T7), .A2(
        top_XOR_T22_U1_xorInst_n9), .ZN(top_XOR_T22_U1_xorInst_n12) );
  INV_X1 top_XOR_T22_U1_xorInst_U1 ( .A(top_T21), .ZN(
        top_XOR_T22_U1_xorInst_n9) );
  AND2_X1 top_XOR_T22_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_189), .A2(
        top_new_AGEMA_signal_180), .ZN(top_XOR_T22_U1_w[0]) );
  AND2_X1 top_XOR_T22_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_190), .A2(
        top_new_AGEMA_signal_179), .ZN(top_XOR_T22_U1_w[1]) );
  AND2_X1 top_XOR_T22_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_190), .A2(
        top_new_AGEMA_signal_180), .ZN(top_XOR_T22_U1_w[2]) );
  AND2_X1 top_XOR_T22_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_189), .A2(
        top_new_AGEMA_signal_179), .ZN(top_XOR_T22_U1_w[3]) );
  OR2_X1 top_XOR_T22_U1_orInst1_U1 ( .A1(top_XOR_T22_U1_w[0]), .A2(
        top_XOR_T22_U1_w[1]), .ZN(top_new_AGEMA_signal_203) );
  OR2_X1 top_XOR_T22_U1_orInst2_U1 ( .A1(top_XOR_T22_U1_w[2]), .A2(
        top_XOR_T22_U1_w[3]), .ZN(top_new_AGEMA_signal_204) );
  OR2_X1 top_XOR_T23_U1_xorInst_U5 ( .A1(top_XOR_T23_U1_xorInst_n12), .A2(
        top_XOR_T23_U1_xorInst_n11), .ZN(top_T23) );
  INV_X1 top_XOR_T23_U1_xorInst_U4 ( .A(top_XOR_T23_U1_xorInst_n10), .ZN(
        top_XOR_T23_U1_xorInst_n11) );
  OR2_X1 top_XOR_T23_U1_xorInst_U3 ( .A1(top_XOR_T23_U1_xorInst_n9), .A2(
        top_T2), .ZN(top_XOR_T23_U1_xorInst_n10) );
  AND2_X1 top_XOR_T23_U1_xorInst_U2 ( .A1(top_T2), .A2(
        top_XOR_T23_U1_xorInst_n9), .ZN(top_XOR_T23_U1_xorInst_n12) );
  INV_X1 top_XOR_T23_U1_xorInst_U1 ( .A(top_T22), .ZN(
        top_XOR_T23_U1_xorInst_n9) );
  AND2_X1 top_XOR_T23_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_203), .A2(
        top_new_AGEMA_signal_164), .ZN(top_XOR_T23_U1_w[0]) );
  AND2_X1 top_XOR_T23_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_204), .A2(
        top_new_AGEMA_signal_163), .ZN(top_XOR_T23_U1_w[1]) );
  AND2_X1 top_XOR_T23_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_204), .A2(
        top_new_AGEMA_signal_164), .ZN(top_XOR_T23_U1_w[2]) );
  AND2_X1 top_XOR_T23_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_203), .A2(
        top_new_AGEMA_signal_163), .ZN(top_XOR_T23_U1_w[3]) );
  OR2_X1 top_XOR_T23_U1_orInst1_U1 ( .A1(top_XOR_T23_U1_w[0]), .A2(
        top_XOR_T23_U1_w[1]), .ZN(top_new_AGEMA_signal_217) );
  OR2_X1 top_XOR_T23_U1_orInst2_U1 ( .A1(top_XOR_T23_U1_w[2]), .A2(
        top_XOR_T23_U1_w[3]), .ZN(top_new_AGEMA_signal_218) );
  OR2_X1 top_XOR_T24_U1_xorInst_U5 ( .A1(top_XOR_T24_U1_xorInst_n12), .A2(
        top_XOR_T24_U1_xorInst_n11), .ZN(top_T24) );
  INV_X1 top_XOR_T24_U1_xorInst_U4 ( .A(top_XOR_T24_U1_xorInst_n10), .ZN(
        top_XOR_T24_U1_xorInst_n11) );
  OR2_X1 top_XOR_T24_U1_xorInst_U3 ( .A1(top_XOR_T24_U1_xorInst_n9), .A2(
        top_T2), .ZN(top_XOR_T24_U1_xorInst_n10) );
  AND2_X1 top_XOR_T24_U1_xorInst_U2 ( .A1(top_T2), .A2(
        top_XOR_T24_U1_xorInst_n9), .ZN(top_XOR_T24_U1_xorInst_n12) );
  INV_X1 top_XOR_T24_U1_xorInst_U1 ( .A(top_T10), .ZN(
        top_XOR_T24_U1_xorInst_n9) );
  AND2_X1 top_XOR_T24_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_209), .A2(
        top_new_AGEMA_signal_164), .ZN(top_XOR_T24_U1_w[0]) );
  AND2_X1 top_XOR_T24_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_210), .A2(
        top_new_AGEMA_signal_163), .ZN(top_XOR_T24_U1_w[1]) );
  AND2_X1 top_XOR_T24_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_210), .A2(
        top_new_AGEMA_signal_164), .ZN(top_XOR_T24_U1_w[2]) );
  AND2_X1 top_XOR_T24_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_209), .A2(
        top_new_AGEMA_signal_163), .ZN(top_XOR_T24_U1_w[3]) );
  OR2_X1 top_XOR_T24_U1_orInst1_U1 ( .A1(top_XOR_T24_U1_w[0]), .A2(
        top_XOR_T24_U1_w[1]), .ZN(top_new_AGEMA_signal_233) );
  OR2_X1 top_XOR_T24_U1_orInst2_U1 ( .A1(top_XOR_T24_U1_w[2]), .A2(
        top_XOR_T24_U1_w[3]), .ZN(top_new_AGEMA_signal_234) );
  OR2_X1 top_XOR_T25_U1_xorInst_U5 ( .A1(top_XOR_T25_U1_xorInst_n12), .A2(
        top_XOR_T25_U1_xorInst_n11), .ZN(top_T25) );
  INV_X1 top_XOR_T25_U1_xorInst_U4 ( .A(top_XOR_T25_U1_xorInst_n10), .ZN(
        top_XOR_T25_U1_xorInst_n11) );
  OR2_X1 top_XOR_T25_U1_xorInst_U3 ( .A1(top_XOR_T25_U1_xorInst_n9), .A2(
        top_T20), .ZN(top_XOR_T25_U1_xorInst_n10) );
  AND2_X1 top_XOR_T25_U1_xorInst_U2 ( .A1(top_T20), .A2(
        top_XOR_T25_U1_xorInst_n9), .ZN(top_XOR_T25_U1_xorInst_n12) );
  INV_X1 top_XOR_T25_U1_xorInst_U1 ( .A(top_T17), .ZN(
        top_XOR_T25_U1_xorInst_n9) );
  AND2_X1 top_XOR_T25_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_213), .A2(
        top_new_AGEMA_signal_216), .ZN(top_XOR_T25_U1_w[0]) );
  AND2_X1 top_XOR_T25_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_214), .A2(
        top_new_AGEMA_signal_215), .ZN(top_XOR_T25_U1_w[1]) );
  AND2_X1 top_XOR_T25_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_214), .A2(
        top_new_AGEMA_signal_216), .ZN(top_XOR_T25_U1_w[2]) );
  AND2_X1 top_XOR_T25_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_213), .A2(
        top_new_AGEMA_signal_215), .ZN(top_XOR_T25_U1_w[3]) );
  OR2_X1 top_XOR_T25_U1_orInst1_U1 ( .A1(top_XOR_T25_U1_w[0]), .A2(
        top_XOR_T25_U1_w[1]), .ZN(top_new_AGEMA_signal_235) );
  OR2_X1 top_XOR_T25_U1_orInst2_U1 ( .A1(top_XOR_T25_U1_w[2]), .A2(
        top_XOR_T25_U1_w[3]), .ZN(top_new_AGEMA_signal_236) );
  OR2_X1 top_XOR_T26_U1_xorInst_U5 ( .A1(top_XOR_T26_U1_xorInst_n12), .A2(
        top_XOR_T26_U1_xorInst_n11), .ZN(top_T26) );
  INV_X1 top_XOR_T26_U1_xorInst_U4 ( .A(top_XOR_T26_U1_xorInst_n10), .ZN(
        top_XOR_T26_U1_xorInst_n11) );
  OR2_X1 top_XOR_T26_U1_xorInst_U3 ( .A1(top_XOR_T26_U1_xorInst_n9), .A2(
        top_T3), .ZN(top_XOR_T26_U1_xorInst_n10) );
  AND2_X1 top_XOR_T26_U1_xorInst_U2 ( .A1(top_T3), .A2(
        top_XOR_T26_U1_xorInst_n9), .ZN(top_XOR_T26_U1_xorInst_n12) );
  INV_X1 top_XOR_T26_U1_xorInst_U1 ( .A(top_T16), .ZN(
        top_XOR_T26_U1_xorInst_n9) );
  AND2_X1 top_XOR_T26_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_199), .A2(
        top_new_AGEMA_signal_168), .ZN(top_XOR_T26_U1_w[0]) );
  AND2_X1 top_XOR_T26_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_200), .A2(
        top_new_AGEMA_signal_167), .ZN(top_XOR_T26_U1_w[1]) );
  AND2_X1 top_XOR_T26_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_200), .A2(
        top_new_AGEMA_signal_168), .ZN(top_XOR_T26_U1_w[2]) );
  AND2_X1 top_XOR_T26_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_199), .A2(
        top_new_AGEMA_signal_167), .ZN(top_XOR_T26_U1_w[3]) );
  OR2_X1 top_XOR_T26_U1_orInst1_U1 ( .A1(top_XOR_T26_U1_w[0]), .A2(
        top_XOR_T26_U1_w[1]), .ZN(top_new_AGEMA_signal_219) );
  OR2_X1 top_XOR_T26_U1_orInst2_U1 ( .A1(top_XOR_T26_U1_w[2]), .A2(
        top_XOR_T26_U1_w[3]), .ZN(top_new_AGEMA_signal_220) );
  OR2_X1 top_XOR_T27_U1_xorInst_U5 ( .A1(top_XOR_T27_U1_xorInst_n12), .A2(
        top_XOR_T27_U1_xorInst_n11), .ZN(top_T27) );
  INV_X1 top_XOR_T27_U1_xorInst_U4 ( .A(top_XOR_T27_U1_xorInst_n10), .ZN(
        top_XOR_T27_U1_xorInst_n11) );
  OR2_X1 top_XOR_T27_U1_xorInst_U3 ( .A1(top_XOR_T27_U1_xorInst_n9), .A2(
        top_T1), .ZN(top_XOR_T27_U1_xorInst_n10) );
  AND2_X1 top_XOR_T27_U1_xorInst_U2 ( .A1(top_T1), .A2(
        top_XOR_T27_U1_xorInst_n9), .ZN(top_XOR_T27_U1_xorInst_n12) );
  INV_X1 top_XOR_T27_U1_xorInst_U1 ( .A(top_T12), .ZN(
        top_XOR_T27_U1_xorInst_n9) );
  AND2_X1 top_XOR_T27_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_183), .A2(
        top_new_AGEMA_signal_160), .ZN(top_XOR_T27_U1_w[0]) );
  AND2_X1 top_XOR_T27_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_184), .A2(
        top_new_AGEMA_signal_159), .ZN(top_XOR_T27_U1_w[1]) );
  AND2_X1 top_XOR_T27_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_184), .A2(
        top_new_AGEMA_signal_160), .ZN(top_XOR_T27_U1_w[2]) );
  AND2_X1 top_XOR_T27_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_183), .A2(
        top_new_AGEMA_signal_159), .ZN(top_XOR_T27_U1_w[3]) );
  OR2_X1 top_XOR_T27_U1_orInst1_U1 ( .A1(top_XOR_T27_U1_w[0]), .A2(
        top_XOR_T27_U1_w[1]), .ZN(top_new_AGEMA_signal_205) );
  OR2_X1 top_XOR_T27_U1_orInst2_U1 ( .A1(top_XOR_T27_U1_w[2]), .A2(
        top_XOR_T27_U1_w[3]), .ZN(top_new_AGEMA_signal_206) );
  INV_X1 top_AND_M1_U1_nonlinearInst_U26 ( .A(top_AND_M1_U1_t[3]), .ZN(
        top_AND_M1_U1_t[7]) );
  OR2_X1 top_AND_M1_U1_nonlinearInst_U25 ( .A1(top_AND_M1_U1_nonlinearInst_n18), .A2(top_AND_M1_U1_nonlinearInst_n17), .ZN(top_AND_M1_U1_t[3]) );
  INV_X1 top_AND_M1_U1_nonlinearInst_U24 ( .A(top_AND_M1_U1_nonlinearInst_n16), 
        .ZN(top_AND_M1_U1_nonlinearInst_n17) );
  OR2_X1 top_AND_M1_U1_nonlinearInst_U23 ( .A1(top_AND_M1_U1_nonlinearInst_n15), .A2(Fresh[0]), .ZN(top_AND_M1_U1_nonlinearInst_n16) );
  AND2_X1 top_AND_M1_U1_nonlinearInst_U22 ( .A1(Fresh[0]), .A2(
        top_AND_M1_U1_nonlinearInst_n15), .ZN(top_AND_M1_U1_nonlinearInst_n18)
         );
  OR2_X1 top_AND_M1_U1_nonlinearInst_U21 ( .A1(top_T13), .A2(top_T6), .ZN(
        top_AND_M1_U1_nonlinearInst_n15) );
  INV_X1 top_AND_M1_U1_nonlinearInst_U20 ( .A(top_AND_M1_U1_t[2]), .ZN(
        top_AND_M1_U1_t[6]) );
  OR2_X1 top_AND_M1_U1_nonlinearInst_U19 ( .A1(top_AND_M1_U1_nonlinearInst_n14), .A2(top_AND_M1_U1_nonlinearInst_n13), .ZN(top_AND_M1_U1_t[2]) );
  INV_X1 top_AND_M1_U1_nonlinearInst_U18 ( .A(top_AND_M1_U1_nonlinearInst_n12), 
        .ZN(top_AND_M1_U1_nonlinearInst_n13) );
  OR2_X1 top_AND_M1_U1_nonlinearInst_U17 ( .A1(top_AND_M1_U1_nonlinearInst_n11), .A2(Fresh[0]), .ZN(top_AND_M1_U1_nonlinearInst_n12) );
  AND2_X1 top_AND_M1_U1_nonlinearInst_U16 ( .A1(Fresh[0]), .A2(
        top_AND_M1_U1_nonlinearInst_n11), .ZN(top_AND_M1_U1_nonlinearInst_n14)
         );
  OR2_X1 top_AND_M1_U1_nonlinearInst_U15 ( .A1(top_AND_M1_U1_nonlinearInst_n10), .A2(top_T13), .ZN(top_AND_M1_U1_nonlinearInst_n11) );
  INV_X1 top_AND_M1_U1_nonlinearInst_U14 ( .A(top_AND_M1_U1_t[1]), .ZN(
        top_AND_M1_U1_t[5]) );
  OR2_X1 top_AND_M1_U1_nonlinearInst_U13 ( .A1(top_AND_M1_U1_nonlinearInst_n9), 
        .A2(top_AND_M1_U1_nonlinearInst_n8), .ZN(top_AND_M1_U1_t[1]) );
  AND2_X1 top_AND_M1_U1_nonlinearInst_U12 ( .A1(top_AND_M1_U1_nonlinearInst_n7), .A2(top_AND_M1_U1_nonlinearInst_n6), .ZN(top_AND_M1_U1_nonlinearInst_n8) );
  INV_X1 top_AND_M1_U1_nonlinearInst_U11 ( .A(top_AND_M1_U1_nonlinearInst_n5), 
        .ZN(top_AND_M1_U1_nonlinearInst_n9) );
  OR2_X1 top_AND_M1_U1_nonlinearInst_U10 ( .A1(top_AND_M1_U1_nonlinearInst_n6), 
        .A2(top_AND_M1_U1_nonlinearInst_n7), .ZN(
        top_AND_M1_U1_nonlinearInst_n5) );
  AND2_X1 top_AND_M1_U1_nonlinearInst_U9 ( .A1(top_T13), .A2(
        top_AND_M1_U1_nonlinearInst_n10), .ZN(top_AND_M1_U1_nonlinearInst_n7)
         );
  INV_X1 top_AND_M1_U1_nonlinearInst_U8 ( .A(top_T6), .ZN(
        top_AND_M1_U1_nonlinearInst_n10) );
  INV_X1 top_AND_M1_U1_nonlinearInst_U7 ( .A(top_AND_M1_U1_t[0]), .ZN(
        top_AND_M1_U1_t[4]) );
  OR2_X1 top_AND_M1_U1_nonlinearInst_U6 ( .A1(top_AND_M1_U1_nonlinearInst_n4), 
        .A2(top_AND_M1_U1_nonlinearInst_n3), .ZN(top_AND_M1_U1_t[0]) );
  AND2_X1 top_AND_M1_U1_nonlinearInst_U5 ( .A1(top_AND_M1_U1_nonlinearInst_n2), 
        .A2(top_AND_M1_U1_nonlinearInst_n6), .ZN(
        top_AND_M1_U1_nonlinearInst_n3) );
  INV_X1 top_AND_M1_U1_nonlinearInst_U4 ( .A(top_AND_M1_U1_nonlinearInst_n1), 
        .ZN(top_AND_M1_U1_nonlinearInst_n4) );
  OR2_X1 top_AND_M1_U1_nonlinearInst_U3 ( .A1(top_AND_M1_U1_nonlinearInst_n6), 
        .A2(top_AND_M1_U1_nonlinearInst_n2), .ZN(
        top_AND_M1_U1_nonlinearInst_n1) );
  AND2_X1 top_AND_M1_U1_nonlinearInst_U2 ( .A1(top_T13), .A2(top_T6), .ZN(
        top_AND_M1_U1_nonlinearInst_n2) );
  INV_X1 top_AND_M1_U1_nonlinearInst_U1 ( .A(Fresh[0]), .ZN(
        top_AND_M1_U1_nonlinearInst_n6) );
  AND2_X1 top_AND_M1_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M1_U1_t[0]), .A2(
        top_AND_M1_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M1_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M1_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M1_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M1_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M1_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M1_U1_t_reg[0]) );
  AND2_X1 top_AND_M1_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M1_U1_t[1]), .A2(
        top_AND_M1_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M1_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M1_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M1_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M1_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M1_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M1_U1_t_reg[1]) );
  AND2_X1 top_AND_M1_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M1_U1_t[2]), .A2(
        top_AND_M1_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M1_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M1_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M1_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M1_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M1_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M1_U1_t_reg[2]) );
  AND2_X1 top_AND_M1_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M1_U1_t[3]), .A2(
        top_AND_M1_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M1_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M1_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M1_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M1_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M1_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M1_U1_t_reg[3]) );
  AND2_X1 top_AND_M1_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M1_U1_t[4]), .A2(
        top_AND_M1_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M1_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M1_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M1_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M1_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M1_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M1_U1_t_reg[4]) );
  AND2_X1 top_AND_M1_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M1_U1_t[5]), .A2(
        top_AND_M1_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M1_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M1_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M1_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M1_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M1_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M1_U1_t_reg[5]) );
  AND2_X1 top_AND_M1_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M1_U1_t[6]), .A2(
        top_AND_M1_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M1_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M1_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M1_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M1_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M1_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M1_U1_t_reg[6]) );
  AND2_X1 top_AND_M1_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M1_U1_t[7]), .A2(
        top_AND_M1_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M1_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M1_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M1_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M1_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M1_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M1_U1_t_reg[7]) );
  AND2_X1 top_AND_M1_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_192), .A2(top_AND_M1_U1_OperationInst_andInst0_n1), .ZN(top_AND_M1_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M1_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_196), .A2(top_AND_M1_U1_t_reg[0]), .ZN(
        top_AND_M1_U1_OperationInst_andInst0_n1) );
  AND2_X1 top_AND_M1_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_191), .A2(top_AND_M1_U1_OperationInst_andInst1_n3), .ZN(top_AND_M1_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M1_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_196), .A2(top_AND_M1_U1_t_reg[1]), .ZN(
        top_AND_M1_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M1_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_192), .A2(top_AND_M1_U1_OperationInst_andInst2_n3), .ZN(top_AND_M1_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M1_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_195), .A2(top_AND_M1_U1_t_reg[2]), .ZN(
        top_AND_M1_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M1_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_191), .A2(top_AND_M1_U1_OperationInst_andInst3_n3), .ZN(top_AND_M1_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M1_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_195), .A2(top_AND_M1_U1_t_reg[3]), .ZN(
        top_AND_M1_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M1_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M1_U1_OperationInst_q[1]), .A2(
        top_AND_M1_U1_OperationInst_orInst1_n2), .ZN(top_new_AGEMA_signal_221)
         );
  OR2_X1 top_AND_M1_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M1_U1_OperationInst_q[0]), .A2(
        top_AND_M1_U1_OperationInst_orInst1_n1), .ZN(
        top_AND_M1_U1_OperationInst_orInst1_n2) );
  OR2_X1 top_AND_M1_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M1_U1_OperationInst_q[3]), .A2(
        top_AND_M1_U1_OperationInst_q[2]), .ZN(
        top_AND_M1_U1_OperationInst_orInst1_n1) );
  AND2_X1 top_AND_M1_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_192), .A2(top_AND_M1_U1_OperationInst_andInst4_n3), .ZN(top_AND_M1_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M1_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_196), .A2(top_AND_M1_U1_t_reg[4]), .ZN(
        top_AND_M1_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M1_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_191), .A2(top_AND_M1_U1_OperationInst_andInst5_n3), .ZN(top_AND_M1_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M1_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_196), .A2(top_AND_M1_U1_t_reg[5]), .ZN(
        top_AND_M1_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M1_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_192), .A2(top_AND_M1_U1_OperationInst_andInst6_n3), .ZN(top_AND_M1_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M1_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_195), .A2(top_AND_M1_U1_t_reg[6]), .ZN(
        top_AND_M1_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M1_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_191), .A2(top_AND_M1_U1_OperationInst_andInst7_n3), .ZN(top_AND_M1_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M1_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_195), .A2(top_AND_M1_U1_t_reg[7]), .ZN(
        top_AND_M1_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M1_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M1_U1_OperationInst_q[5]), .A2(
        top_AND_M1_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_222)
         );
  OR2_X1 top_AND_M1_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M1_U1_OperationInst_q[4]), .A2(
        top_AND_M1_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M1_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M1_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M1_U1_OperationInst_q[7]), .A2(
        top_AND_M1_U1_OperationInst_q[6]), .ZN(
        top_AND_M1_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M2_U1_nonlinearInst_U26 ( .A(top_AND_M2_U1_t[3]), .ZN(
        top_AND_M2_U1_t[7]) );
  OR2_X1 top_AND_M2_U1_nonlinearInst_U25 ( .A1(top_AND_M2_U1_nonlinearInst_n64), .A2(top_AND_M2_U1_nonlinearInst_n63), .ZN(top_AND_M2_U1_t[3]) );
  INV_X1 top_AND_M2_U1_nonlinearInst_U24 ( .A(top_AND_M2_U1_nonlinearInst_n62), 
        .ZN(top_AND_M2_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M2_U1_nonlinearInst_U23 ( .A1(top_AND_M2_U1_nonlinearInst_n61), .A2(Fresh[1]), .ZN(top_AND_M2_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M2_U1_nonlinearInst_U22 ( .A1(Fresh[1]), .A2(
        top_AND_M2_U1_nonlinearInst_n61), .ZN(top_AND_M2_U1_nonlinearInst_n64)
         );
  OR2_X1 top_AND_M2_U1_nonlinearInst_U21 ( .A1(top_T23), .A2(top_T8), .ZN(
        top_AND_M2_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M2_U1_nonlinearInst_U20 ( .A(top_AND_M2_U1_t[2]), .ZN(
        top_AND_M2_U1_t[6]) );
  OR2_X1 top_AND_M2_U1_nonlinearInst_U19 ( .A1(top_AND_M2_U1_nonlinearInst_n60), .A2(top_AND_M2_U1_nonlinearInst_n59), .ZN(top_AND_M2_U1_t[2]) );
  INV_X1 top_AND_M2_U1_nonlinearInst_U18 ( .A(top_AND_M2_U1_nonlinearInst_n58), 
        .ZN(top_AND_M2_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M2_U1_nonlinearInst_U17 ( .A1(top_AND_M2_U1_nonlinearInst_n57), .A2(Fresh[1]), .ZN(top_AND_M2_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M2_U1_nonlinearInst_U16 ( .A1(Fresh[1]), .A2(
        top_AND_M2_U1_nonlinearInst_n57), .ZN(top_AND_M2_U1_nonlinearInst_n60)
         );
  OR2_X1 top_AND_M2_U1_nonlinearInst_U15 ( .A1(top_AND_M2_U1_nonlinearInst_n56), .A2(top_T23), .ZN(top_AND_M2_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M2_U1_nonlinearInst_U14 ( .A(top_AND_M2_U1_t[1]), .ZN(
        top_AND_M2_U1_t[5]) );
  OR2_X1 top_AND_M2_U1_nonlinearInst_U13 ( .A1(top_AND_M2_U1_nonlinearInst_n55), .A2(top_AND_M2_U1_nonlinearInst_n54), .ZN(top_AND_M2_U1_t[1]) );
  AND2_X1 top_AND_M2_U1_nonlinearInst_U12 ( .A1(
        top_AND_M2_U1_nonlinearInst_n53), .A2(top_AND_M2_U1_nonlinearInst_n52), 
        .ZN(top_AND_M2_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M2_U1_nonlinearInst_U11 ( .A(top_AND_M2_U1_nonlinearInst_n51), 
        .ZN(top_AND_M2_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M2_U1_nonlinearInst_U10 ( .A1(top_AND_M2_U1_nonlinearInst_n52), .A2(top_AND_M2_U1_nonlinearInst_n53), .ZN(top_AND_M2_U1_nonlinearInst_n51)
         );
  AND2_X1 top_AND_M2_U1_nonlinearInst_U9 ( .A1(top_T23), .A2(
        top_AND_M2_U1_nonlinearInst_n56), .ZN(top_AND_M2_U1_nonlinearInst_n53)
         );
  INV_X1 top_AND_M2_U1_nonlinearInst_U8 ( .A(top_T8), .ZN(
        top_AND_M2_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M2_U1_nonlinearInst_U7 ( .A(top_AND_M2_U1_t[0]), .ZN(
        top_AND_M2_U1_t[4]) );
  OR2_X1 top_AND_M2_U1_nonlinearInst_U6 ( .A1(top_AND_M2_U1_nonlinearInst_n50), 
        .A2(top_AND_M2_U1_nonlinearInst_n49), .ZN(top_AND_M2_U1_t[0]) );
  AND2_X1 top_AND_M2_U1_nonlinearInst_U5 ( .A1(top_AND_M2_U1_nonlinearInst_n48), .A2(top_AND_M2_U1_nonlinearInst_n52), .ZN(top_AND_M2_U1_nonlinearInst_n49)
         );
  INV_X1 top_AND_M2_U1_nonlinearInst_U4 ( .A(top_AND_M2_U1_nonlinearInst_n47), 
        .ZN(top_AND_M2_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M2_U1_nonlinearInst_U3 ( .A1(top_AND_M2_U1_nonlinearInst_n52), 
        .A2(top_AND_M2_U1_nonlinearInst_n48), .ZN(
        top_AND_M2_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M2_U1_nonlinearInst_U2 ( .A1(top_T23), .A2(top_T8), .ZN(
        top_AND_M2_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M2_U1_nonlinearInst_U1 ( .A(Fresh[1]), .ZN(
        top_AND_M2_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M2_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M2_U1_t[0]), .A2(
        top_AND_M2_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M2_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M2_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M2_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M2_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M2_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M2_U1_t_reg[0]) );
  AND2_X1 top_AND_M2_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M2_U1_t[1]), .A2(
        top_AND_M2_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M2_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M2_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M2_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M2_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M2_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M2_U1_t_reg[1]) );
  AND2_X1 top_AND_M2_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M2_U1_t[2]), .A2(
        top_AND_M2_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M2_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M2_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M2_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M2_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M2_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M2_U1_t_reg[2]) );
  AND2_X1 top_AND_M2_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M2_U1_t[3]), .A2(
        top_AND_M2_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M2_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M2_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M2_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M2_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M2_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M2_U1_t_reg[3]) );
  AND2_X1 top_AND_M2_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M2_U1_t[4]), .A2(
        top_AND_M2_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M2_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M2_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M2_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M2_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M2_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M2_U1_t_reg[4]) );
  AND2_X1 top_AND_M2_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M2_U1_t[5]), .A2(
        top_AND_M2_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M2_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M2_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M2_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M2_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M2_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M2_U1_t_reg[5]) );
  AND2_X1 top_AND_M2_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M2_U1_t[6]), .A2(
        top_AND_M2_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M2_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M2_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M2_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M2_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M2_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M2_U1_t_reg[6]) );
  AND2_X1 top_AND_M2_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M2_U1_t[7]), .A2(
        top_AND_M2_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M2_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M2_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M2_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M2_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M2_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M2_U1_t_reg[7]) );
  AND2_X1 top_AND_M2_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_208), .A2(top_AND_M2_U1_OperationInst_andInst0_n3), .ZN(top_AND_M2_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M2_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_218), .A2(top_AND_M2_U1_t_reg[0]), .ZN(
        top_AND_M2_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M2_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_207), .A2(top_AND_M2_U1_OperationInst_andInst1_n3), .ZN(top_AND_M2_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M2_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_218), .A2(top_AND_M2_U1_t_reg[1]), .ZN(
        top_AND_M2_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M2_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_208), .A2(top_AND_M2_U1_OperationInst_andInst2_n3), .ZN(top_AND_M2_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M2_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_217), .A2(top_AND_M2_U1_t_reg[2]), .ZN(
        top_AND_M2_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M2_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_207), .A2(top_AND_M2_U1_OperationInst_andInst3_n3), .ZN(top_AND_M2_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M2_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_217), .A2(top_AND_M2_U1_t_reg[3]), .ZN(
        top_AND_M2_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M2_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M2_U1_OperationInst_q[1]), .A2(
        top_AND_M2_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_237)
         );
  OR2_X1 top_AND_M2_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M2_U1_OperationInst_q[0]), .A2(
        top_AND_M2_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M2_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M2_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M2_U1_OperationInst_q[3]), .A2(
        top_AND_M2_U1_OperationInst_q[2]), .ZN(
        top_AND_M2_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M2_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_208), .A2(top_AND_M2_U1_OperationInst_andInst4_n3), .ZN(top_AND_M2_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M2_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_218), .A2(top_AND_M2_U1_t_reg[4]), .ZN(
        top_AND_M2_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M2_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_207), .A2(top_AND_M2_U1_OperationInst_andInst5_n3), .ZN(top_AND_M2_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M2_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_218), .A2(top_AND_M2_U1_t_reg[5]), .ZN(
        top_AND_M2_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M2_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_208), .A2(top_AND_M2_U1_OperationInst_andInst6_n3), .ZN(top_AND_M2_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M2_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_217), .A2(top_AND_M2_U1_t_reg[6]), .ZN(
        top_AND_M2_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M2_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_207), .A2(top_AND_M2_U1_OperationInst_andInst7_n3), .ZN(top_AND_M2_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M2_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_217), .A2(top_AND_M2_U1_t_reg[7]), .ZN(
        top_AND_M2_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M2_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M2_U1_OperationInst_q[5]), .A2(
        top_AND_M2_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_238)
         );
  OR2_X1 top_AND_M2_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M2_U1_OperationInst_q[4]), .A2(
        top_AND_M2_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M2_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M2_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M2_U1_OperationInst_q[7]), .A2(
        top_AND_M2_U1_OperationInst_q[6]), .ZN(
        top_AND_M2_U1_OperationInst_orInst2_n5) );
  OR2_X1 top_XOR_M3_U1_xorInst_U5 ( .A1(top_XOR_M3_U1_xorInst_n12), .A2(
        top_XOR_M3_U1_xorInst_n11), .ZN(top_M3) );
  INV_X1 top_XOR_M3_U1_xorInst_U4 ( .A(top_XOR_M3_U1_xorInst_n10), .ZN(
        top_XOR_M3_U1_xorInst_n11) );
  OR2_X1 top_XOR_M3_U1_xorInst_U3 ( .A1(top_XOR_M3_U1_xorInst_n9), .A2(top_T14), .ZN(top_XOR_M3_U1_xorInst_n10) );
  AND2_X1 top_XOR_M3_U1_xorInst_U2 ( .A1(top_T14), .A2(
        top_XOR_M3_U1_xorInst_n9), .ZN(top_XOR_M3_U1_xorInst_n12) );
  INV_X1 top_XOR_M3_U1_xorInst_U1 ( .A(Fresh[0]), .ZN(top_XOR_M3_U1_xorInst_n9) );
  AND2_X1 top_XOR_M3_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_221), .A2(
        top_new_AGEMA_signal_212), .ZN(top_XOR_M3_U1_w[0]) );
  AND2_X1 top_XOR_M3_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_222), .A2(
        top_new_AGEMA_signal_211), .ZN(top_XOR_M3_U1_w[1]) );
  AND2_X1 top_XOR_M3_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_222), .A2(
        top_new_AGEMA_signal_212), .ZN(top_XOR_M3_U1_w[2]) );
  AND2_X1 top_XOR_M3_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_221), .A2(
        top_new_AGEMA_signal_211), .ZN(top_XOR_M3_U1_w[3]) );
  OR2_X1 top_XOR_M3_U1_orInst1_U1 ( .A1(top_XOR_M3_U1_w[0]), .A2(
        top_XOR_M3_U1_w[1]), .ZN(top_new_AGEMA_signal_239) );
  OR2_X1 top_XOR_M3_U1_orInst2_U1 ( .A1(top_XOR_M3_U1_w[2]), .A2(
        top_XOR_M3_U1_w[3]), .ZN(top_new_AGEMA_signal_240) );
  INV_X1 top_AND_M4_U1_nonlinearInst_U26 ( .A(top_AND_M4_U1_t[3]), .ZN(
        top_AND_M4_U1_t[7]) );
  OR2_X1 top_AND_M4_U1_nonlinearInst_U25 ( .A1(top_AND_M4_U1_nonlinearInst_n64), .A2(top_AND_M4_U1_nonlinearInst_n63), .ZN(top_AND_M4_U1_t[3]) );
  INV_X1 top_AND_M4_U1_nonlinearInst_U24 ( .A(top_AND_M4_U1_nonlinearInst_n62), 
        .ZN(top_AND_M4_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M4_U1_nonlinearInst_U23 ( .A1(top_AND_M4_U1_nonlinearInst_n61), .A2(Fresh[2]), .ZN(top_AND_M4_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M4_U1_nonlinearInst_U22 ( .A1(Fresh[2]), .A2(
        top_AND_M4_U1_nonlinearInst_n61), .ZN(top_AND_M4_U1_nonlinearInst_n64)
         );
  OR2_X1 top_AND_M4_U1_nonlinearInst_U21 ( .A1(top_T19), .A2(X_s0[0]), .ZN(
        top_AND_M4_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M4_U1_nonlinearInst_U20 ( .A(top_AND_M4_U1_t[2]), .ZN(
        top_AND_M4_U1_t[6]) );
  OR2_X1 top_AND_M4_U1_nonlinearInst_U19 ( .A1(top_AND_M4_U1_nonlinearInst_n60), .A2(top_AND_M4_U1_nonlinearInst_n59), .ZN(top_AND_M4_U1_t[2]) );
  INV_X1 top_AND_M4_U1_nonlinearInst_U18 ( .A(top_AND_M4_U1_nonlinearInst_n58), 
        .ZN(top_AND_M4_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M4_U1_nonlinearInst_U17 ( .A1(top_AND_M4_U1_nonlinearInst_n57), .A2(Fresh[2]), .ZN(top_AND_M4_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M4_U1_nonlinearInst_U16 ( .A1(Fresh[2]), .A2(
        top_AND_M4_U1_nonlinearInst_n57), .ZN(top_AND_M4_U1_nonlinearInst_n60)
         );
  OR2_X1 top_AND_M4_U1_nonlinearInst_U15 ( .A1(top_AND_M4_U1_nonlinearInst_n56), .A2(top_T19), .ZN(top_AND_M4_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M4_U1_nonlinearInst_U14 ( .A(top_AND_M4_U1_t[1]), .ZN(
        top_AND_M4_U1_t[5]) );
  OR2_X1 top_AND_M4_U1_nonlinearInst_U13 ( .A1(top_AND_M4_U1_nonlinearInst_n55), .A2(top_AND_M4_U1_nonlinearInst_n54), .ZN(top_AND_M4_U1_t[1]) );
  AND2_X1 top_AND_M4_U1_nonlinearInst_U12 ( .A1(
        top_AND_M4_U1_nonlinearInst_n53), .A2(top_AND_M4_U1_nonlinearInst_n52), 
        .ZN(top_AND_M4_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M4_U1_nonlinearInst_U11 ( .A(top_AND_M4_U1_nonlinearInst_n51), 
        .ZN(top_AND_M4_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M4_U1_nonlinearInst_U10 ( .A1(top_AND_M4_U1_nonlinearInst_n52), .A2(top_AND_M4_U1_nonlinearInst_n53), .ZN(top_AND_M4_U1_nonlinearInst_n51)
         );
  AND2_X1 top_AND_M4_U1_nonlinearInst_U9 ( .A1(top_T19), .A2(
        top_AND_M4_U1_nonlinearInst_n56), .ZN(top_AND_M4_U1_nonlinearInst_n53)
         );
  INV_X1 top_AND_M4_U1_nonlinearInst_U8 ( .A(X_s0[0]), .ZN(
        top_AND_M4_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M4_U1_nonlinearInst_U7 ( .A(top_AND_M4_U1_t[0]), .ZN(
        top_AND_M4_U1_t[4]) );
  OR2_X1 top_AND_M4_U1_nonlinearInst_U6 ( .A1(top_AND_M4_U1_nonlinearInst_n50), 
        .A2(top_AND_M4_U1_nonlinearInst_n49), .ZN(top_AND_M4_U1_t[0]) );
  AND2_X1 top_AND_M4_U1_nonlinearInst_U5 ( .A1(top_AND_M4_U1_nonlinearInst_n48), .A2(top_AND_M4_U1_nonlinearInst_n52), .ZN(top_AND_M4_U1_nonlinearInst_n49)
         );
  INV_X1 top_AND_M4_U1_nonlinearInst_U4 ( .A(top_AND_M4_U1_nonlinearInst_n47), 
        .ZN(top_AND_M4_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M4_U1_nonlinearInst_U3 ( .A1(top_AND_M4_U1_nonlinearInst_n52), 
        .A2(top_AND_M4_U1_nonlinearInst_n48), .ZN(
        top_AND_M4_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M4_U1_nonlinearInst_U2 ( .A1(top_T19), .A2(X_s0[0]), .ZN(
        top_AND_M4_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M4_U1_nonlinearInst_U1 ( .A(Fresh[2]), .ZN(
        top_AND_M4_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M4_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M4_U1_t[0]), .A2(
        top_AND_M4_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M4_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M4_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M4_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M4_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M4_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M4_U1_t_reg[0]) );
  AND2_X1 top_AND_M4_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M4_U1_t[1]), .A2(
        top_AND_M4_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M4_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M4_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M4_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M4_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M4_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M4_U1_t_reg[1]) );
  AND2_X1 top_AND_M4_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M4_U1_t[2]), .A2(
        top_AND_M4_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M4_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M4_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M4_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M4_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M4_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M4_U1_t_reg[2]) );
  AND2_X1 top_AND_M4_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M4_U1_t[3]), .A2(
        top_AND_M4_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M4_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M4_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M4_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M4_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M4_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M4_U1_t_reg[3]) );
  AND2_X1 top_AND_M4_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M4_U1_t[4]), .A2(
        top_AND_M4_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M4_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M4_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M4_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M4_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M4_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M4_U1_t_reg[4]) );
  AND2_X1 top_AND_M4_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M4_U1_t[5]), .A2(
        top_AND_M4_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M4_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M4_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M4_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M4_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M4_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M4_U1_t_reg[5]) );
  AND2_X1 top_AND_M4_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M4_U1_t[6]), .A2(
        top_AND_M4_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M4_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M4_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M4_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M4_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M4_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M4_U1_t_reg[6]) );
  AND2_X1 top_AND_M4_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M4_U1_t[7]), .A2(
        top_AND_M4_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M4_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M4_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M4_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M4_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M4_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M4_U1_t_reg[7]) );
  AND2_X1 top_AND_M4_U1_OperationInst_andInst0_U2 ( .A1(X_s1_bar[0]), .A2(
        top_AND_M4_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M4_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M4_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_202), .A2(top_AND_M4_U1_t_reg[0]), .ZN(
        top_AND_M4_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M4_U1_OperationInst_andInst1_U2 ( .A1(X_s1[0]), .A2(
        top_AND_M4_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M4_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M4_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_202), .A2(top_AND_M4_U1_t_reg[1]), .ZN(
        top_AND_M4_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M4_U1_OperationInst_andInst2_U2 ( .A1(X_s1_bar[0]), .A2(
        top_AND_M4_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M4_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M4_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_201), .A2(top_AND_M4_U1_t_reg[2]), .ZN(
        top_AND_M4_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M4_U1_OperationInst_andInst3_U2 ( .A1(X_s1[0]), .A2(
        top_AND_M4_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M4_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M4_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_201), .A2(top_AND_M4_U1_t_reg[3]), .ZN(
        top_AND_M4_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M4_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M4_U1_OperationInst_q[1]), .A2(
        top_AND_M4_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_223)
         );
  OR2_X1 top_AND_M4_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M4_U1_OperationInst_q[0]), .A2(
        top_AND_M4_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M4_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M4_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M4_U1_OperationInst_q[3]), .A2(
        top_AND_M4_U1_OperationInst_q[2]), .ZN(
        top_AND_M4_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M4_U1_OperationInst_andInst4_U2 ( .A1(X_s1_bar[0]), .A2(
        top_AND_M4_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M4_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M4_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_202), .A2(top_AND_M4_U1_t_reg[4]), .ZN(
        top_AND_M4_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M4_U1_OperationInst_andInst5_U2 ( .A1(X_s1[0]), .A2(
        top_AND_M4_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M4_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M4_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_202), .A2(top_AND_M4_U1_t_reg[5]), .ZN(
        top_AND_M4_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M4_U1_OperationInst_andInst6_U2 ( .A1(X_s1_bar[0]), .A2(
        top_AND_M4_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M4_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M4_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_201), .A2(top_AND_M4_U1_t_reg[6]), .ZN(
        top_AND_M4_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M4_U1_OperationInst_andInst7_U2 ( .A1(X_s1[0]), .A2(
        top_AND_M4_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M4_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M4_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_201), .A2(top_AND_M4_U1_t_reg[7]), .ZN(
        top_AND_M4_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M4_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M4_U1_OperationInst_q[5]), .A2(
        top_AND_M4_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_224)
         );
  OR2_X1 top_AND_M4_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M4_U1_OperationInst_q[4]), .A2(
        top_AND_M4_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M4_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M4_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M4_U1_OperationInst_q[7]), .A2(
        top_AND_M4_U1_OperationInst_q[6]), .ZN(
        top_AND_M4_U1_OperationInst_orInst2_n5) );
  OR2_X1 top_XOR_M5_U1_xorInst_U5 ( .A1(top_XOR_M5_U1_xorInst_n12), .A2(
        top_XOR_M5_U1_xorInst_n11), .ZN(top_M5) );
  INV_X1 top_XOR_M5_U1_xorInst_U4 ( .A(top_XOR_M5_U1_xorInst_n10), .ZN(
        top_XOR_M5_U1_xorInst_n11) );
  OR2_X1 top_XOR_M5_U1_xorInst_U3 ( .A1(top_XOR_M5_U1_xorInst_n9), .A2(
        Fresh[2]), .ZN(top_XOR_M5_U1_xorInst_n10) );
  AND2_X1 top_XOR_M5_U1_xorInst_U2 ( .A1(Fresh[2]), .A2(
        top_XOR_M5_U1_xorInst_n9), .ZN(top_XOR_M5_U1_xorInst_n12) );
  INV_X1 top_XOR_M5_U1_xorInst_U1 ( .A(Fresh[0]), .ZN(top_XOR_M5_U1_xorInst_n9) );
  AND2_X1 top_XOR_M5_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_221), .A2(
        top_new_AGEMA_signal_224), .ZN(top_XOR_M5_U1_w[0]) );
  AND2_X1 top_XOR_M5_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_222), .A2(
        top_new_AGEMA_signal_223), .ZN(top_XOR_M5_U1_w[1]) );
  AND2_X1 top_XOR_M5_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_222), .A2(
        top_new_AGEMA_signal_224), .ZN(top_XOR_M5_U1_w[2]) );
  AND2_X1 top_XOR_M5_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_221), .A2(
        top_new_AGEMA_signal_223), .ZN(top_XOR_M5_U1_w[3]) );
  OR2_X1 top_XOR_M5_U1_orInst1_U1 ( .A1(top_XOR_M5_U1_w[0]), .A2(
        top_XOR_M5_U1_w[1]), .ZN(top_new_AGEMA_signal_241) );
  OR2_X1 top_XOR_M5_U1_orInst2_U1 ( .A1(top_XOR_M5_U1_w[2]), .A2(
        top_XOR_M5_U1_w[3]), .ZN(top_new_AGEMA_signal_242) );
  INV_X1 top_AND_M6_U1_nonlinearInst_U26 ( .A(top_AND_M6_U1_t[3]), .ZN(
        top_AND_M6_U1_t[7]) );
  OR2_X1 top_AND_M6_U1_nonlinearInst_U25 ( .A1(top_AND_M6_U1_nonlinearInst_n64), .A2(top_AND_M6_U1_nonlinearInst_n63), .ZN(top_AND_M6_U1_t[3]) );
  INV_X1 top_AND_M6_U1_nonlinearInst_U24 ( .A(top_AND_M6_U1_nonlinearInst_n62), 
        .ZN(top_AND_M6_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M6_U1_nonlinearInst_U23 ( .A1(top_AND_M6_U1_nonlinearInst_n61), .A2(Fresh[3]), .ZN(top_AND_M6_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M6_U1_nonlinearInst_U22 ( .A1(Fresh[3]), .A2(
        top_AND_M6_U1_nonlinearInst_n61), .ZN(top_AND_M6_U1_nonlinearInst_n64)
         );
  OR2_X1 top_AND_M6_U1_nonlinearInst_U21 ( .A1(top_T3), .A2(top_T16), .ZN(
        top_AND_M6_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M6_U1_nonlinearInst_U20 ( .A(top_AND_M6_U1_t[2]), .ZN(
        top_AND_M6_U1_t[6]) );
  OR2_X1 top_AND_M6_U1_nonlinearInst_U19 ( .A1(top_AND_M6_U1_nonlinearInst_n60), .A2(top_AND_M6_U1_nonlinearInst_n59), .ZN(top_AND_M6_U1_t[2]) );
  INV_X1 top_AND_M6_U1_nonlinearInst_U18 ( .A(top_AND_M6_U1_nonlinearInst_n58), 
        .ZN(top_AND_M6_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M6_U1_nonlinearInst_U17 ( .A1(top_AND_M6_U1_nonlinearInst_n57), .A2(Fresh[3]), .ZN(top_AND_M6_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M6_U1_nonlinearInst_U16 ( .A1(Fresh[3]), .A2(
        top_AND_M6_U1_nonlinearInst_n57), .ZN(top_AND_M6_U1_nonlinearInst_n60)
         );
  OR2_X1 top_AND_M6_U1_nonlinearInst_U15 ( .A1(top_AND_M6_U1_nonlinearInst_n56), .A2(top_T3), .ZN(top_AND_M6_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M6_U1_nonlinearInst_U14 ( .A(top_AND_M6_U1_t[1]), .ZN(
        top_AND_M6_U1_t[5]) );
  OR2_X1 top_AND_M6_U1_nonlinearInst_U13 ( .A1(top_AND_M6_U1_nonlinearInst_n55), .A2(top_AND_M6_U1_nonlinearInst_n54), .ZN(top_AND_M6_U1_t[1]) );
  AND2_X1 top_AND_M6_U1_nonlinearInst_U12 ( .A1(
        top_AND_M6_U1_nonlinearInst_n53), .A2(top_AND_M6_U1_nonlinearInst_n52), 
        .ZN(top_AND_M6_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M6_U1_nonlinearInst_U11 ( .A(top_AND_M6_U1_nonlinearInst_n51), 
        .ZN(top_AND_M6_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M6_U1_nonlinearInst_U10 ( .A1(top_AND_M6_U1_nonlinearInst_n52), .A2(top_AND_M6_U1_nonlinearInst_n53), .ZN(top_AND_M6_U1_nonlinearInst_n51)
         );
  AND2_X1 top_AND_M6_U1_nonlinearInst_U9 ( .A1(top_T3), .A2(
        top_AND_M6_U1_nonlinearInst_n56), .ZN(top_AND_M6_U1_nonlinearInst_n53)
         );
  INV_X1 top_AND_M6_U1_nonlinearInst_U8 ( .A(top_T16), .ZN(
        top_AND_M6_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M6_U1_nonlinearInst_U7 ( .A(top_AND_M6_U1_t[0]), .ZN(
        top_AND_M6_U1_t[4]) );
  OR2_X1 top_AND_M6_U1_nonlinearInst_U6 ( .A1(top_AND_M6_U1_nonlinearInst_n50), 
        .A2(top_AND_M6_U1_nonlinearInst_n49), .ZN(top_AND_M6_U1_t[0]) );
  AND2_X1 top_AND_M6_U1_nonlinearInst_U5 ( .A1(top_AND_M6_U1_nonlinearInst_n48), .A2(top_AND_M6_U1_nonlinearInst_n52), .ZN(top_AND_M6_U1_nonlinearInst_n49)
         );
  INV_X1 top_AND_M6_U1_nonlinearInst_U4 ( .A(top_AND_M6_U1_nonlinearInst_n47), 
        .ZN(top_AND_M6_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M6_U1_nonlinearInst_U3 ( .A1(top_AND_M6_U1_nonlinearInst_n52), 
        .A2(top_AND_M6_U1_nonlinearInst_n48), .ZN(
        top_AND_M6_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M6_U1_nonlinearInst_U2 ( .A1(top_T3), .A2(top_T16), .ZN(
        top_AND_M6_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M6_U1_nonlinearInst_U1 ( .A(Fresh[3]), .ZN(
        top_AND_M6_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M6_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M6_U1_t[0]), .A2(
        top_AND_M6_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M6_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M6_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M6_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M6_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M6_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M6_U1_t_reg[0]) );
  AND2_X1 top_AND_M6_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M6_U1_t[1]), .A2(
        top_AND_M6_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M6_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M6_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M6_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M6_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M6_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M6_U1_t_reg[1]) );
  AND2_X1 top_AND_M6_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M6_U1_t[2]), .A2(
        top_AND_M6_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M6_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M6_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M6_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M6_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M6_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M6_U1_t_reg[2]) );
  AND2_X1 top_AND_M6_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M6_U1_t[3]), .A2(
        top_AND_M6_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M6_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M6_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M6_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M6_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M6_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M6_U1_t_reg[3]) );
  AND2_X1 top_AND_M6_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M6_U1_t[4]), .A2(
        top_AND_M6_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M6_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M6_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M6_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M6_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M6_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M6_U1_t_reg[4]) );
  AND2_X1 top_AND_M6_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M6_U1_t[5]), .A2(
        top_AND_M6_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M6_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M6_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M6_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M6_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M6_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M6_U1_t_reg[5]) );
  AND2_X1 top_AND_M6_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M6_U1_t[6]), .A2(
        top_AND_M6_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M6_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M6_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M6_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M6_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M6_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M6_U1_t_reg[6]) );
  AND2_X1 top_AND_M6_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M6_U1_t[7]), .A2(
        top_AND_M6_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M6_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M6_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M6_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M6_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M6_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M6_U1_t_reg[7]) );
  AND2_X1 top_AND_M6_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_200), .A2(top_AND_M6_U1_OperationInst_andInst0_n3), .ZN(top_AND_M6_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M6_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_168), .A2(top_AND_M6_U1_t_reg[0]), .ZN(
        top_AND_M6_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M6_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_199), .A2(top_AND_M6_U1_OperationInst_andInst1_n3), .ZN(top_AND_M6_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M6_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_168), .A2(top_AND_M6_U1_t_reg[1]), .ZN(
        top_AND_M6_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M6_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_200), .A2(top_AND_M6_U1_OperationInst_andInst2_n3), .ZN(top_AND_M6_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M6_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_167), .A2(top_AND_M6_U1_t_reg[2]), .ZN(
        top_AND_M6_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M6_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_199), .A2(top_AND_M6_U1_OperationInst_andInst3_n3), .ZN(top_AND_M6_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M6_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_167), .A2(top_AND_M6_U1_t_reg[3]), .ZN(
        top_AND_M6_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M6_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M6_U1_OperationInst_q[1]), .A2(
        top_AND_M6_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_225)
         );
  OR2_X1 top_AND_M6_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M6_U1_OperationInst_q[0]), .A2(
        top_AND_M6_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M6_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M6_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M6_U1_OperationInst_q[3]), .A2(
        top_AND_M6_U1_OperationInst_q[2]), .ZN(
        top_AND_M6_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M6_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_200), .A2(top_AND_M6_U1_OperationInst_andInst4_n3), .ZN(top_AND_M6_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M6_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_168), .A2(top_AND_M6_U1_t_reg[4]), .ZN(
        top_AND_M6_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M6_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_199), .A2(top_AND_M6_U1_OperationInst_andInst5_n3), .ZN(top_AND_M6_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M6_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_168), .A2(top_AND_M6_U1_t_reg[5]), .ZN(
        top_AND_M6_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M6_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_200), .A2(top_AND_M6_U1_OperationInst_andInst6_n3), .ZN(top_AND_M6_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M6_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_167), .A2(top_AND_M6_U1_t_reg[6]), .ZN(
        top_AND_M6_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M6_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_199), .A2(top_AND_M6_U1_OperationInst_andInst7_n3), .ZN(top_AND_M6_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M6_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_167), .A2(top_AND_M6_U1_t_reg[7]), .ZN(
        top_AND_M6_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M6_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M6_U1_OperationInst_q[5]), .A2(
        top_AND_M6_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_226)
         );
  OR2_X1 top_AND_M6_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M6_U1_OperationInst_q[4]), .A2(
        top_AND_M6_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M6_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M6_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M6_U1_OperationInst_q[7]), .A2(
        top_AND_M6_U1_OperationInst_q[6]), .ZN(
        top_AND_M6_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M7_U1_nonlinearInst_U26 ( .A(top_AND_M7_U1_t[3]), .ZN(
        top_AND_M7_U1_t[7]) );
  OR2_X1 top_AND_M7_U1_nonlinearInst_U25 ( .A1(top_AND_M7_U1_nonlinearInst_n64), .A2(top_AND_M7_U1_nonlinearInst_n63), .ZN(top_AND_M7_U1_t[3]) );
  INV_X1 top_AND_M7_U1_nonlinearInst_U24 ( .A(top_AND_M7_U1_nonlinearInst_n62), 
        .ZN(top_AND_M7_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M7_U1_nonlinearInst_U23 ( .A1(top_AND_M7_U1_nonlinearInst_n61), .A2(Fresh[4]), .ZN(top_AND_M7_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M7_U1_nonlinearInst_U22 ( .A1(Fresh[4]), .A2(
        top_AND_M7_U1_nonlinearInst_n61), .ZN(top_AND_M7_U1_nonlinearInst_n64)
         );
  OR2_X1 top_AND_M7_U1_nonlinearInst_U21 ( .A1(top_T22), .A2(top_T9), .ZN(
        top_AND_M7_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M7_U1_nonlinearInst_U20 ( .A(top_AND_M7_U1_t[2]), .ZN(
        top_AND_M7_U1_t[6]) );
  OR2_X1 top_AND_M7_U1_nonlinearInst_U19 ( .A1(top_AND_M7_U1_nonlinearInst_n60), .A2(top_AND_M7_U1_nonlinearInst_n59), .ZN(top_AND_M7_U1_t[2]) );
  INV_X1 top_AND_M7_U1_nonlinearInst_U18 ( .A(top_AND_M7_U1_nonlinearInst_n58), 
        .ZN(top_AND_M7_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M7_U1_nonlinearInst_U17 ( .A1(top_AND_M7_U1_nonlinearInst_n57), .A2(Fresh[4]), .ZN(top_AND_M7_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M7_U1_nonlinearInst_U16 ( .A1(Fresh[4]), .A2(
        top_AND_M7_U1_nonlinearInst_n57), .ZN(top_AND_M7_U1_nonlinearInst_n60)
         );
  OR2_X1 top_AND_M7_U1_nonlinearInst_U15 ( .A1(top_AND_M7_U1_nonlinearInst_n56), .A2(top_T22), .ZN(top_AND_M7_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M7_U1_nonlinearInst_U14 ( .A(top_AND_M7_U1_t[1]), .ZN(
        top_AND_M7_U1_t[5]) );
  OR2_X1 top_AND_M7_U1_nonlinearInst_U13 ( .A1(top_AND_M7_U1_nonlinearInst_n55), .A2(top_AND_M7_U1_nonlinearInst_n54), .ZN(top_AND_M7_U1_t[1]) );
  AND2_X1 top_AND_M7_U1_nonlinearInst_U12 ( .A1(
        top_AND_M7_U1_nonlinearInst_n53), .A2(top_AND_M7_U1_nonlinearInst_n52), 
        .ZN(top_AND_M7_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M7_U1_nonlinearInst_U11 ( .A(top_AND_M7_U1_nonlinearInst_n51), 
        .ZN(top_AND_M7_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M7_U1_nonlinearInst_U10 ( .A1(top_AND_M7_U1_nonlinearInst_n52), .A2(top_AND_M7_U1_nonlinearInst_n53), .ZN(top_AND_M7_U1_nonlinearInst_n51)
         );
  AND2_X1 top_AND_M7_U1_nonlinearInst_U9 ( .A1(top_T22), .A2(
        top_AND_M7_U1_nonlinearInst_n56), .ZN(top_AND_M7_U1_nonlinearInst_n53)
         );
  INV_X1 top_AND_M7_U1_nonlinearInst_U8 ( .A(top_T9), .ZN(
        top_AND_M7_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M7_U1_nonlinearInst_U7 ( .A(top_AND_M7_U1_t[0]), .ZN(
        top_AND_M7_U1_t[4]) );
  OR2_X1 top_AND_M7_U1_nonlinearInst_U6 ( .A1(top_AND_M7_U1_nonlinearInst_n50), 
        .A2(top_AND_M7_U1_nonlinearInst_n49), .ZN(top_AND_M7_U1_t[0]) );
  AND2_X1 top_AND_M7_U1_nonlinearInst_U5 ( .A1(top_AND_M7_U1_nonlinearInst_n48), .A2(top_AND_M7_U1_nonlinearInst_n52), .ZN(top_AND_M7_U1_nonlinearInst_n49)
         );
  INV_X1 top_AND_M7_U1_nonlinearInst_U4 ( .A(top_AND_M7_U1_nonlinearInst_n47), 
        .ZN(top_AND_M7_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M7_U1_nonlinearInst_U3 ( .A1(top_AND_M7_U1_nonlinearInst_n52), 
        .A2(top_AND_M7_U1_nonlinearInst_n48), .ZN(
        top_AND_M7_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M7_U1_nonlinearInst_U2 ( .A1(top_T22), .A2(top_T9), .ZN(
        top_AND_M7_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M7_U1_nonlinearInst_U1 ( .A(Fresh[4]), .ZN(
        top_AND_M7_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M7_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M7_U1_t[0]), .A2(
        top_AND_M7_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M7_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M7_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M7_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M7_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M7_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M7_U1_t_reg[0]) );
  AND2_X1 top_AND_M7_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M7_U1_t[1]), .A2(
        top_AND_M7_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M7_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M7_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M7_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M7_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M7_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M7_U1_t_reg[1]) );
  AND2_X1 top_AND_M7_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M7_U1_t[2]), .A2(
        top_AND_M7_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M7_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M7_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M7_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M7_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M7_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M7_U1_t_reg[2]) );
  AND2_X1 top_AND_M7_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M7_U1_t[3]), .A2(
        top_AND_M7_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M7_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M7_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M7_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M7_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M7_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M7_U1_t_reg[3]) );
  AND2_X1 top_AND_M7_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M7_U1_t[4]), .A2(
        top_AND_M7_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M7_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M7_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M7_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M7_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M7_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M7_U1_t_reg[4]) );
  AND2_X1 top_AND_M7_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M7_U1_t[5]), .A2(
        top_AND_M7_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M7_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M7_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M7_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M7_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M7_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M7_U1_t_reg[5]) );
  AND2_X1 top_AND_M7_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M7_U1_t[6]), .A2(
        top_AND_M7_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M7_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M7_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M7_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M7_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M7_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M7_U1_t_reg[6]) );
  AND2_X1 top_AND_M7_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M7_U1_t[7]), .A2(
        top_AND_M7_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M7_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M7_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M7_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M7_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M7_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M7_U1_t_reg[7]) );
  AND2_X1 top_AND_M7_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_194), .A2(top_AND_M7_U1_OperationInst_andInst0_n3), .ZN(top_AND_M7_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M7_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_204), .A2(top_AND_M7_U1_t_reg[0]), .ZN(
        top_AND_M7_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M7_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_193), .A2(top_AND_M7_U1_OperationInst_andInst1_n3), .ZN(top_AND_M7_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M7_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_204), .A2(top_AND_M7_U1_t_reg[1]), .ZN(
        top_AND_M7_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M7_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_194), .A2(top_AND_M7_U1_OperationInst_andInst2_n3), .ZN(top_AND_M7_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M7_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_203), .A2(top_AND_M7_U1_t_reg[2]), .ZN(
        top_AND_M7_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M7_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_193), .A2(top_AND_M7_U1_OperationInst_andInst3_n3), .ZN(top_AND_M7_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M7_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_203), .A2(top_AND_M7_U1_t_reg[3]), .ZN(
        top_AND_M7_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M7_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M7_U1_OperationInst_q[1]), .A2(
        top_AND_M7_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_227)
         );
  OR2_X1 top_AND_M7_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M7_U1_OperationInst_q[0]), .A2(
        top_AND_M7_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M7_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M7_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M7_U1_OperationInst_q[3]), .A2(
        top_AND_M7_U1_OperationInst_q[2]), .ZN(
        top_AND_M7_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M7_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_194), .A2(top_AND_M7_U1_OperationInst_andInst4_n3), .ZN(top_AND_M7_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M7_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_204), .A2(top_AND_M7_U1_t_reg[4]), .ZN(
        top_AND_M7_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M7_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_193), .A2(top_AND_M7_U1_OperationInst_andInst5_n3), .ZN(top_AND_M7_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M7_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_204), .A2(top_AND_M7_U1_t_reg[5]), .ZN(
        top_AND_M7_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M7_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_194), .A2(top_AND_M7_U1_OperationInst_andInst6_n3), .ZN(top_AND_M7_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M7_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_203), .A2(top_AND_M7_U1_t_reg[6]), .ZN(
        top_AND_M7_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M7_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_193), .A2(top_AND_M7_U1_OperationInst_andInst7_n3), .ZN(top_AND_M7_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M7_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_203), .A2(top_AND_M7_U1_t_reg[7]), .ZN(
        top_AND_M7_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M7_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M7_U1_OperationInst_q[5]), .A2(
        top_AND_M7_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_228)
         );
  OR2_X1 top_AND_M7_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M7_U1_OperationInst_q[4]), .A2(
        top_AND_M7_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M7_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M7_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M7_U1_OperationInst_q[7]), .A2(
        top_AND_M7_U1_OperationInst_q[6]), .ZN(
        top_AND_M7_U1_OperationInst_orInst2_n5) );
  OR2_X1 top_XOR_M8_U1_xorInst_U5 ( .A1(top_XOR_M8_U1_xorInst_n12), .A2(
        top_XOR_M8_U1_xorInst_n11), .ZN(top_M8) );
  INV_X1 top_XOR_M8_U1_xorInst_U4 ( .A(top_XOR_M8_U1_xorInst_n10), .ZN(
        top_XOR_M8_U1_xorInst_n11) );
  OR2_X1 top_XOR_M8_U1_xorInst_U3 ( .A1(top_XOR_M8_U1_xorInst_n9), .A2(top_T26), .ZN(top_XOR_M8_U1_xorInst_n10) );
  AND2_X1 top_XOR_M8_U1_xorInst_U2 ( .A1(top_T26), .A2(
        top_XOR_M8_U1_xorInst_n9), .ZN(top_XOR_M8_U1_xorInst_n12) );
  INV_X1 top_XOR_M8_U1_xorInst_U1 ( .A(Fresh[3]), .ZN(top_XOR_M8_U1_xorInst_n9) );
  AND2_X1 top_XOR_M8_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_225), .A2(
        top_new_AGEMA_signal_220), .ZN(top_XOR_M8_U1_w[0]) );
  AND2_X1 top_XOR_M8_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_226), .A2(
        top_new_AGEMA_signal_219), .ZN(top_XOR_M8_U1_w[1]) );
  AND2_X1 top_XOR_M8_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_226), .A2(
        top_new_AGEMA_signal_220), .ZN(top_XOR_M8_U1_w[2]) );
  AND2_X1 top_XOR_M8_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_225), .A2(
        top_new_AGEMA_signal_219), .ZN(top_XOR_M8_U1_w[3]) );
  OR2_X1 top_XOR_M8_U1_orInst1_U1 ( .A1(top_XOR_M8_U1_w[0]), .A2(
        top_XOR_M8_U1_w[1]), .ZN(top_new_AGEMA_signal_243) );
  OR2_X1 top_XOR_M8_U1_orInst2_U1 ( .A1(top_XOR_M8_U1_w[2]), .A2(
        top_XOR_M8_U1_w[3]), .ZN(top_new_AGEMA_signal_244) );
  INV_X1 top_AND_M9_U1_nonlinearInst_U26 ( .A(top_AND_M9_U1_t[3]), .ZN(
        top_AND_M9_U1_t[7]) );
  OR2_X1 top_AND_M9_U1_nonlinearInst_U25 ( .A1(top_AND_M9_U1_nonlinearInst_n64), .A2(top_AND_M9_U1_nonlinearInst_n63), .ZN(top_AND_M9_U1_t[3]) );
  INV_X1 top_AND_M9_U1_nonlinearInst_U24 ( .A(top_AND_M9_U1_nonlinearInst_n62), 
        .ZN(top_AND_M9_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M9_U1_nonlinearInst_U23 ( .A1(top_AND_M9_U1_nonlinearInst_n61), .A2(Fresh[5]), .ZN(top_AND_M9_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M9_U1_nonlinearInst_U22 ( .A1(Fresh[5]), .A2(
        top_AND_M9_U1_nonlinearInst_n61), .ZN(top_AND_M9_U1_nonlinearInst_n64)
         );
  OR2_X1 top_AND_M9_U1_nonlinearInst_U21 ( .A1(top_T20), .A2(top_T17), .ZN(
        top_AND_M9_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M9_U1_nonlinearInst_U20 ( .A(top_AND_M9_U1_t[2]), .ZN(
        top_AND_M9_U1_t[6]) );
  OR2_X1 top_AND_M9_U1_nonlinearInst_U19 ( .A1(top_AND_M9_U1_nonlinearInst_n60), .A2(top_AND_M9_U1_nonlinearInst_n59), .ZN(top_AND_M9_U1_t[2]) );
  INV_X1 top_AND_M9_U1_nonlinearInst_U18 ( .A(top_AND_M9_U1_nonlinearInst_n58), 
        .ZN(top_AND_M9_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M9_U1_nonlinearInst_U17 ( .A1(top_AND_M9_U1_nonlinearInst_n57), .A2(Fresh[5]), .ZN(top_AND_M9_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M9_U1_nonlinearInst_U16 ( .A1(Fresh[5]), .A2(
        top_AND_M9_U1_nonlinearInst_n57), .ZN(top_AND_M9_U1_nonlinearInst_n60)
         );
  OR2_X1 top_AND_M9_U1_nonlinearInst_U15 ( .A1(top_AND_M9_U1_nonlinearInst_n56), .A2(top_T20), .ZN(top_AND_M9_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M9_U1_nonlinearInst_U14 ( .A(top_AND_M9_U1_t[1]), .ZN(
        top_AND_M9_U1_t[5]) );
  OR2_X1 top_AND_M9_U1_nonlinearInst_U13 ( .A1(top_AND_M9_U1_nonlinearInst_n55), .A2(top_AND_M9_U1_nonlinearInst_n54), .ZN(top_AND_M9_U1_t[1]) );
  AND2_X1 top_AND_M9_U1_nonlinearInst_U12 ( .A1(
        top_AND_M9_U1_nonlinearInst_n53), .A2(top_AND_M9_U1_nonlinearInst_n52), 
        .ZN(top_AND_M9_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M9_U1_nonlinearInst_U11 ( .A(top_AND_M9_U1_nonlinearInst_n51), 
        .ZN(top_AND_M9_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M9_U1_nonlinearInst_U10 ( .A1(top_AND_M9_U1_nonlinearInst_n52), .A2(top_AND_M9_U1_nonlinearInst_n53), .ZN(top_AND_M9_U1_nonlinearInst_n51)
         );
  AND2_X1 top_AND_M9_U1_nonlinearInst_U9 ( .A1(top_T20), .A2(
        top_AND_M9_U1_nonlinearInst_n56), .ZN(top_AND_M9_U1_nonlinearInst_n53)
         );
  INV_X1 top_AND_M9_U1_nonlinearInst_U8 ( .A(top_T17), .ZN(
        top_AND_M9_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M9_U1_nonlinearInst_U7 ( .A(top_AND_M9_U1_t[0]), .ZN(
        top_AND_M9_U1_t[4]) );
  OR2_X1 top_AND_M9_U1_nonlinearInst_U6 ( .A1(top_AND_M9_U1_nonlinearInst_n50), 
        .A2(top_AND_M9_U1_nonlinearInst_n49), .ZN(top_AND_M9_U1_t[0]) );
  AND2_X1 top_AND_M9_U1_nonlinearInst_U5 ( .A1(top_AND_M9_U1_nonlinearInst_n48), .A2(top_AND_M9_U1_nonlinearInst_n52), .ZN(top_AND_M9_U1_nonlinearInst_n49)
         );
  INV_X1 top_AND_M9_U1_nonlinearInst_U4 ( .A(top_AND_M9_U1_nonlinearInst_n47), 
        .ZN(top_AND_M9_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M9_U1_nonlinearInst_U3 ( .A1(top_AND_M9_U1_nonlinearInst_n52), 
        .A2(top_AND_M9_U1_nonlinearInst_n48), .ZN(
        top_AND_M9_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M9_U1_nonlinearInst_U2 ( .A1(top_T20), .A2(top_T17), .ZN(
        top_AND_M9_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M9_U1_nonlinearInst_U1 ( .A(Fresh[5]), .ZN(
        top_AND_M9_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M9_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M9_U1_t[0]), .A2(
        top_AND_M9_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M9_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M9_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M9_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M9_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M9_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M9_U1_t_reg[0]) );
  AND2_X1 top_AND_M9_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M9_U1_t[1]), .A2(
        top_AND_M9_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M9_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M9_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M9_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M9_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M9_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M9_U1_t_reg[1]) );
  AND2_X1 top_AND_M9_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M9_U1_t[2]), .A2(
        top_AND_M9_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M9_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M9_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M9_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M9_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M9_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M9_U1_t_reg[2]) );
  AND2_X1 top_AND_M9_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M9_U1_t[3]), .A2(
        top_AND_M9_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M9_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M9_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M9_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M9_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M9_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M9_U1_t_reg[3]) );
  AND2_X1 top_AND_M9_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M9_U1_t[4]), .A2(
        top_AND_M9_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M9_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M9_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M9_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M9_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M9_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M9_U1_t_reg[4]) );
  AND2_X1 top_AND_M9_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M9_U1_t[5]), .A2(
        top_AND_M9_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M9_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M9_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M9_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M9_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M9_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M9_U1_t_reg[5]) );
  AND2_X1 top_AND_M9_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M9_U1_t[6]), .A2(
        top_AND_M9_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M9_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M9_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M9_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M9_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M9_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M9_U1_t_reg[6]) );
  AND2_X1 top_AND_M9_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M9_U1_t[7]), .A2(
        top_AND_M9_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M9_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M9_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M9_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M9_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M9_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M9_U1_t_reg[7]) );
  AND2_X1 top_AND_M9_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_214), .A2(top_AND_M9_U1_OperationInst_andInst0_n3), .ZN(top_AND_M9_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M9_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_216), .A2(top_AND_M9_U1_t_reg[0]), .ZN(
        top_AND_M9_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M9_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_213), .A2(top_AND_M9_U1_OperationInst_andInst1_n3), .ZN(top_AND_M9_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M9_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_216), .A2(top_AND_M9_U1_t_reg[1]), .ZN(
        top_AND_M9_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M9_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_214), .A2(top_AND_M9_U1_OperationInst_andInst2_n3), .ZN(top_AND_M9_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M9_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_215), .A2(top_AND_M9_U1_t_reg[2]), .ZN(
        top_AND_M9_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M9_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_213), .A2(top_AND_M9_U1_OperationInst_andInst3_n3), .ZN(top_AND_M9_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M9_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_215), .A2(top_AND_M9_U1_t_reg[3]), .ZN(
        top_AND_M9_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M9_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M9_U1_OperationInst_q[1]), .A2(
        top_AND_M9_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_245)
         );
  OR2_X1 top_AND_M9_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M9_U1_OperationInst_q[0]), .A2(
        top_AND_M9_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M9_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M9_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M9_U1_OperationInst_q[3]), .A2(
        top_AND_M9_U1_OperationInst_q[2]), .ZN(
        top_AND_M9_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M9_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_214), .A2(top_AND_M9_U1_OperationInst_andInst4_n3), .ZN(top_AND_M9_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M9_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_216), .A2(top_AND_M9_U1_t_reg[4]), .ZN(
        top_AND_M9_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M9_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_213), .A2(top_AND_M9_U1_OperationInst_andInst5_n3), .ZN(top_AND_M9_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M9_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_216), .A2(top_AND_M9_U1_t_reg[5]), .ZN(
        top_AND_M9_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M9_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_214), .A2(top_AND_M9_U1_OperationInst_andInst6_n3), .ZN(top_AND_M9_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M9_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_215), .A2(top_AND_M9_U1_t_reg[6]), .ZN(
        top_AND_M9_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M9_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_213), .A2(top_AND_M9_U1_OperationInst_andInst7_n3), .ZN(top_AND_M9_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M9_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_215), .A2(top_AND_M9_U1_t_reg[7]), .ZN(
        top_AND_M9_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M9_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M9_U1_OperationInst_q[5]), .A2(
        top_AND_M9_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_246)
         );
  OR2_X1 top_AND_M9_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M9_U1_OperationInst_q[4]), .A2(
        top_AND_M9_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M9_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M9_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M9_U1_OperationInst_q[7]), .A2(
        top_AND_M9_U1_OperationInst_q[6]), .ZN(
        top_AND_M9_U1_OperationInst_orInst2_n5) );
  OR2_X1 top_XOR_M10_U1_xorInst_U5 ( .A1(top_XOR_M10_U1_xorInst_n12), .A2(
        top_XOR_M10_U1_xorInst_n11), .ZN(top_M10) );
  INV_X1 top_XOR_M10_U1_xorInst_U4 ( .A(top_XOR_M10_U1_xorInst_n10), .ZN(
        top_XOR_M10_U1_xorInst_n11) );
  OR2_X1 top_XOR_M10_U1_xorInst_U3 ( .A1(top_XOR_M10_U1_xorInst_n9), .A2(
        Fresh[5]), .ZN(top_XOR_M10_U1_xorInst_n10) );
  AND2_X1 top_XOR_M10_U1_xorInst_U2 ( .A1(Fresh[5]), .A2(
        top_XOR_M10_U1_xorInst_n9), .ZN(top_XOR_M10_U1_xorInst_n12) );
  INV_X1 top_XOR_M10_U1_xorInst_U1 ( .A(Fresh[3]), .ZN(
        top_XOR_M10_U1_xorInst_n9) );
  AND2_X1 top_XOR_M10_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_225), .A2(
        top_new_AGEMA_signal_246), .ZN(top_XOR_M10_U1_w[0]) );
  AND2_X1 top_XOR_M10_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_226), .A2(
        top_new_AGEMA_signal_245), .ZN(top_XOR_M10_U1_w[1]) );
  AND2_X1 top_XOR_M10_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_226), .A2(
        top_new_AGEMA_signal_246), .ZN(top_XOR_M10_U1_w[2]) );
  AND2_X1 top_XOR_M10_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_225), .A2(
        top_new_AGEMA_signal_245), .ZN(top_XOR_M10_U1_w[3]) );
  OR2_X1 top_XOR_M10_U1_orInst1_U1 ( .A1(top_XOR_M10_U1_w[0]), .A2(
        top_XOR_M10_U1_w[1]), .ZN(top_new_AGEMA_signal_251) );
  OR2_X1 top_XOR_M10_U1_orInst2_U1 ( .A1(top_XOR_M10_U1_w[2]), .A2(
        top_XOR_M10_U1_w[3]), .ZN(top_new_AGEMA_signal_252) );
  INV_X1 top_AND_M11_U1_nonlinearInst_U26 ( .A(top_AND_M11_U1_t[3]), .ZN(
        top_AND_M11_U1_t[7]) );
  OR2_X1 top_AND_M11_U1_nonlinearInst_U25 ( .A1(
        top_AND_M11_U1_nonlinearInst_n64), .A2(
        top_AND_M11_U1_nonlinearInst_n63), .ZN(top_AND_M11_U1_t[3]) );
  INV_X1 top_AND_M11_U1_nonlinearInst_U24 ( .A(
        top_AND_M11_U1_nonlinearInst_n62), .ZN(
        top_AND_M11_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M11_U1_nonlinearInst_U23 ( .A1(
        top_AND_M11_U1_nonlinearInst_n61), .A2(Fresh[6]), .ZN(
        top_AND_M11_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M11_U1_nonlinearInst_U22 ( .A1(Fresh[6]), .A2(
        top_AND_M11_U1_nonlinearInst_n61), .ZN(
        top_AND_M11_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M11_U1_nonlinearInst_U21 ( .A1(top_T1), .A2(top_T15), .ZN(
        top_AND_M11_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M11_U1_nonlinearInst_U20 ( .A(top_AND_M11_U1_t[2]), .ZN(
        top_AND_M11_U1_t[6]) );
  OR2_X1 top_AND_M11_U1_nonlinearInst_U19 ( .A1(
        top_AND_M11_U1_nonlinearInst_n60), .A2(
        top_AND_M11_U1_nonlinearInst_n59), .ZN(top_AND_M11_U1_t[2]) );
  INV_X1 top_AND_M11_U1_nonlinearInst_U18 ( .A(
        top_AND_M11_U1_nonlinearInst_n58), .ZN(
        top_AND_M11_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M11_U1_nonlinearInst_U17 ( .A1(
        top_AND_M11_U1_nonlinearInst_n57), .A2(Fresh[6]), .ZN(
        top_AND_M11_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M11_U1_nonlinearInst_U16 ( .A1(Fresh[6]), .A2(
        top_AND_M11_U1_nonlinearInst_n57), .ZN(
        top_AND_M11_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M11_U1_nonlinearInst_U15 ( .A1(
        top_AND_M11_U1_nonlinearInst_n56), .A2(top_T1), .ZN(
        top_AND_M11_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M11_U1_nonlinearInst_U14 ( .A(top_AND_M11_U1_t[1]), .ZN(
        top_AND_M11_U1_t[5]) );
  OR2_X1 top_AND_M11_U1_nonlinearInst_U13 ( .A1(
        top_AND_M11_U1_nonlinearInst_n55), .A2(
        top_AND_M11_U1_nonlinearInst_n54), .ZN(top_AND_M11_U1_t[1]) );
  AND2_X1 top_AND_M11_U1_nonlinearInst_U12 ( .A1(
        top_AND_M11_U1_nonlinearInst_n53), .A2(
        top_AND_M11_U1_nonlinearInst_n52), .ZN(
        top_AND_M11_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M11_U1_nonlinearInst_U11 ( .A(
        top_AND_M11_U1_nonlinearInst_n51), .ZN(
        top_AND_M11_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M11_U1_nonlinearInst_U10 ( .A1(
        top_AND_M11_U1_nonlinearInst_n52), .A2(
        top_AND_M11_U1_nonlinearInst_n53), .ZN(
        top_AND_M11_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M11_U1_nonlinearInst_U9 ( .A1(top_T1), .A2(
        top_AND_M11_U1_nonlinearInst_n56), .ZN(
        top_AND_M11_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M11_U1_nonlinearInst_U8 ( .A(top_T15), .ZN(
        top_AND_M11_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M11_U1_nonlinearInst_U7 ( .A(top_AND_M11_U1_t[0]), .ZN(
        top_AND_M11_U1_t[4]) );
  OR2_X1 top_AND_M11_U1_nonlinearInst_U6 ( .A1(
        top_AND_M11_U1_nonlinearInst_n50), .A2(
        top_AND_M11_U1_nonlinearInst_n49), .ZN(top_AND_M11_U1_t[0]) );
  AND2_X1 top_AND_M11_U1_nonlinearInst_U5 ( .A1(
        top_AND_M11_U1_nonlinearInst_n48), .A2(
        top_AND_M11_U1_nonlinearInst_n52), .ZN(
        top_AND_M11_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M11_U1_nonlinearInst_U4 ( .A(top_AND_M11_U1_nonlinearInst_n47), .ZN(top_AND_M11_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M11_U1_nonlinearInst_U3 ( .A1(
        top_AND_M11_U1_nonlinearInst_n52), .A2(
        top_AND_M11_U1_nonlinearInst_n48), .ZN(
        top_AND_M11_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M11_U1_nonlinearInst_U2 ( .A1(top_T1), .A2(top_T15), .ZN(
        top_AND_M11_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M11_U1_nonlinearInst_U1 ( .A(Fresh[6]), .ZN(
        top_AND_M11_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M11_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M11_U1_t[0]), .A2(
        top_AND_M11_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M11_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M11_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M11_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M11_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M11_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M11_U1_t_reg[0]) );
  AND2_X1 top_AND_M11_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M11_U1_t[1]), .A2(
        top_AND_M11_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M11_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M11_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M11_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M11_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M11_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M11_U1_t_reg[1]) );
  AND2_X1 top_AND_M11_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M11_U1_t[2]), .A2(
        top_AND_M11_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M11_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M11_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M11_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M11_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M11_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M11_U1_t_reg[2]) );
  AND2_X1 top_AND_M11_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M11_U1_t[3]), .A2(
        top_AND_M11_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M11_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M11_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M11_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M11_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M11_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M11_U1_t_reg[3]) );
  AND2_X1 top_AND_M11_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M11_U1_t[4]), .A2(
        top_AND_M11_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M11_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M11_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M11_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M11_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M11_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M11_U1_t_reg[4]) );
  AND2_X1 top_AND_M11_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M11_U1_t[5]), .A2(
        top_AND_M11_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M11_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M11_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M11_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M11_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M11_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M11_U1_t_reg[5]) );
  AND2_X1 top_AND_M11_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M11_U1_t[6]), .A2(
        top_AND_M11_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M11_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M11_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M11_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M11_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M11_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M11_U1_t_reg[6]) );
  AND2_X1 top_AND_M11_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M11_U1_t[7]), .A2(
        top_AND_M11_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M11_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M11_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M11_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M11_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M11_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M11_U1_t_reg[7]) );
  AND2_X1 top_AND_M11_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_198), .A2(
        top_AND_M11_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M11_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M11_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_160), .A2(top_AND_M11_U1_t_reg[0]), .ZN(
        top_AND_M11_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M11_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_197), .A2(
        top_AND_M11_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M11_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M11_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_160), .A2(top_AND_M11_U1_t_reg[1]), .ZN(
        top_AND_M11_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M11_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_198), .A2(
        top_AND_M11_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M11_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M11_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_159), .A2(top_AND_M11_U1_t_reg[2]), .ZN(
        top_AND_M11_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M11_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_197), .A2(
        top_AND_M11_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M11_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M11_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_159), .A2(top_AND_M11_U1_t_reg[3]), .ZN(
        top_AND_M11_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M11_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M11_U1_OperationInst_q[1]), .A2(
        top_AND_M11_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_229) );
  OR2_X1 top_AND_M11_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M11_U1_OperationInst_q[0]), .A2(
        top_AND_M11_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M11_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M11_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M11_U1_OperationInst_q[3]), .A2(
        top_AND_M11_U1_OperationInst_q[2]), .ZN(
        top_AND_M11_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M11_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_198), .A2(
        top_AND_M11_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M11_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M11_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_160), .A2(top_AND_M11_U1_t_reg[4]), .ZN(
        top_AND_M11_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M11_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_197), .A2(
        top_AND_M11_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M11_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M11_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_160), .A2(top_AND_M11_U1_t_reg[5]), .ZN(
        top_AND_M11_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M11_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_198), .A2(
        top_AND_M11_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M11_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M11_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_159), .A2(top_AND_M11_U1_t_reg[6]), .ZN(
        top_AND_M11_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M11_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_197), .A2(
        top_AND_M11_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M11_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M11_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_159), .A2(top_AND_M11_U1_t_reg[7]), .ZN(
        top_AND_M11_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M11_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M11_U1_OperationInst_q[5]), .A2(
        top_AND_M11_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_230) );
  OR2_X1 top_AND_M11_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M11_U1_OperationInst_q[4]), .A2(
        top_AND_M11_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M11_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M11_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M11_U1_OperationInst_q[7]), .A2(
        top_AND_M11_U1_OperationInst_q[6]), .ZN(
        top_AND_M11_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M12_U1_nonlinearInst_U26 ( .A(top_AND_M12_U1_t[3]), .ZN(
        top_AND_M12_U1_t[7]) );
  OR2_X1 top_AND_M12_U1_nonlinearInst_U25 ( .A1(
        top_AND_M12_U1_nonlinearInst_n64), .A2(
        top_AND_M12_U1_nonlinearInst_n63), .ZN(top_AND_M12_U1_t[3]) );
  INV_X1 top_AND_M12_U1_nonlinearInst_U24 ( .A(
        top_AND_M12_U1_nonlinearInst_n62), .ZN(
        top_AND_M12_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M12_U1_nonlinearInst_U23 ( .A1(
        top_AND_M12_U1_nonlinearInst_n61), .A2(Fresh[7]), .ZN(
        top_AND_M12_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M12_U1_nonlinearInst_U22 ( .A1(Fresh[7]), .A2(
        top_AND_M12_U1_nonlinearInst_n61), .ZN(
        top_AND_M12_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M12_U1_nonlinearInst_U21 ( .A1(top_T4), .A2(top_T27), .ZN(
        top_AND_M12_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M12_U1_nonlinearInst_U20 ( .A(top_AND_M12_U1_t[2]), .ZN(
        top_AND_M12_U1_t[6]) );
  OR2_X1 top_AND_M12_U1_nonlinearInst_U19 ( .A1(
        top_AND_M12_U1_nonlinearInst_n60), .A2(
        top_AND_M12_U1_nonlinearInst_n59), .ZN(top_AND_M12_U1_t[2]) );
  INV_X1 top_AND_M12_U1_nonlinearInst_U18 ( .A(
        top_AND_M12_U1_nonlinearInst_n58), .ZN(
        top_AND_M12_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M12_U1_nonlinearInst_U17 ( .A1(
        top_AND_M12_U1_nonlinearInst_n57), .A2(Fresh[7]), .ZN(
        top_AND_M12_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M12_U1_nonlinearInst_U16 ( .A1(Fresh[7]), .A2(
        top_AND_M12_U1_nonlinearInst_n57), .ZN(
        top_AND_M12_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M12_U1_nonlinearInst_U15 ( .A1(
        top_AND_M12_U1_nonlinearInst_n56), .A2(top_T4), .ZN(
        top_AND_M12_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M12_U1_nonlinearInst_U14 ( .A(top_AND_M12_U1_t[1]), .ZN(
        top_AND_M12_U1_t[5]) );
  OR2_X1 top_AND_M12_U1_nonlinearInst_U13 ( .A1(
        top_AND_M12_U1_nonlinearInst_n55), .A2(
        top_AND_M12_U1_nonlinearInst_n54), .ZN(top_AND_M12_U1_t[1]) );
  AND2_X1 top_AND_M12_U1_nonlinearInst_U12 ( .A1(
        top_AND_M12_U1_nonlinearInst_n53), .A2(
        top_AND_M12_U1_nonlinearInst_n52), .ZN(
        top_AND_M12_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M12_U1_nonlinearInst_U11 ( .A(
        top_AND_M12_U1_nonlinearInst_n51), .ZN(
        top_AND_M12_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M12_U1_nonlinearInst_U10 ( .A1(
        top_AND_M12_U1_nonlinearInst_n52), .A2(
        top_AND_M12_U1_nonlinearInst_n53), .ZN(
        top_AND_M12_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M12_U1_nonlinearInst_U9 ( .A1(top_T4), .A2(
        top_AND_M12_U1_nonlinearInst_n56), .ZN(
        top_AND_M12_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M12_U1_nonlinearInst_U8 ( .A(top_T27), .ZN(
        top_AND_M12_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M12_U1_nonlinearInst_U7 ( .A(top_AND_M12_U1_t[0]), .ZN(
        top_AND_M12_U1_t[4]) );
  OR2_X1 top_AND_M12_U1_nonlinearInst_U6 ( .A1(
        top_AND_M12_U1_nonlinearInst_n50), .A2(
        top_AND_M12_U1_nonlinearInst_n49), .ZN(top_AND_M12_U1_t[0]) );
  AND2_X1 top_AND_M12_U1_nonlinearInst_U5 ( .A1(
        top_AND_M12_U1_nonlinearInst_n48), .A2(
        top_AND_M12_U1_nonlinearInst_n52), .ZN(
        top_AND_M12_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M12_U1_nonlinearInst_U4 ( .A(top_AND_M12_U1_nonlinearInst_n47), .ZN(top_AND_M12_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M12_U1_nonlinearInst_U3 ( .A1(
        top_AND_M12_U1_nonlinearInst_n52), .A2(
        top_AND_M12_U1_nonlinearInst_n48), .ZN(
        top_AND_M12_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M12_U1_nonlinearInst_U2 ( .A1(top_T4), .A2(top_T27), .ZN(
        top_AND_M12_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M12_U1_nonlinearInst_U1 ( .A(Fresh[7]), .ZN(
        top_AND_M12_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M12_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M12_U1_t[0]), .A2(
        top_AND_M12_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M12_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M12_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M12_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M12_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M12_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M12_U1_t_reg[0]) );
  AND2_X1 top_AND_M12_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M12_U1_t[1]), .A2(
        top_AND_M12_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M12_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M12_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M12_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M12_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M12_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M12_U1_t_reg[1]) );
  AND2_X1 top_AND_M12_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M12_U1_t[2]), .A2(
        top_AND_M12_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M12_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M12_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M12_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M12_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M12_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M12_U1_t_reg[2]) );
  AND2_X1 top_AND_M12_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M12_U1_t[3]), .A2(
        top_AND_M12_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M12_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M12_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M12_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M12_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M12_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M12_U1_t_reg[3]) );
  AND2_X1 top_AND_M12_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M12_U1_t[4]), .A2(
        top_AND_M12_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M12_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M12_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M12_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M12_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M12_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M12_U1_t_reg[4]) );
  AND2_X1 top_AND_M12_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M12_U1_t[5]), .A2(
        top_AND_M12_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M12_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M12_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M12_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M12_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M12_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M12_U1_t_reg[5]) );
  AND2_X1 top_AND_M12_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M12_U1_t[6]), .A2(
        top_AND_M12_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M12_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M12_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M12_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M12_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M12_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M12_U1_t_reg[6]) );
  AND2_X1 top_AND_M12_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M12_U1_t[7]), .A2(
        top_AND_M12_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M12_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M12_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M12_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M12_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M12_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M12_U1_t_reg[7]) );
  AND2_X1 top_AND_M12_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_206), .A2(
        top_AND_M12_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M12_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M12_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_170), .A2(top_AND_M12_U1_t_reg[0]), .ZN(
        top_AND_M12_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M12_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_205), .A2(
        top_AND_M12_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M12_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M12_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_170), .A2(top_AND_M12_U1_t_reg[1]), .ZN(
        top_AND_M12_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M12_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_206), .A2(
        top_AND_M12_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M12_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M12_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_169), .A2(top_AND_M12_U1_t_reg[2]), .ZN(
        top_AND_M12_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M12_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_205), .A2(
        top_AND_M12_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M12_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M12_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_169), .A2(top_AND_M12_U1_t_reg[3]), .ZN(
        top_AND_M12_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M12_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M12_U1_OperationInst_q[1]), .A2(
        top_AND_M12_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_231) );
  OR2_X1 top_AND_M12_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M12_U1_OperationInst_q[0]), .A2(
        top_AND_M12_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M12_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M12_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M12_U1_OperationInst_q[3]), .A2(
        top_AND_M12_U1_OperationInst_q[2]), .ZN(
        top_AND_M12_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M12_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_206), .A2(
        top_AND_M12_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M12_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M12_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_170), .A2(top_AND_M12_U1_t_reg[4]), .ZN(
        top_AND_M12_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M12_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_205), .A2(
        top_AND_M12_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M12_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M12_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_170), .A2(top_AND_M12_U1_t_reg[5]), .ZN(
        top_AND_M12_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M12_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_206), .A2(
        top_AND_M12_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M12_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M12_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_169), .A2(top_AND_M12_U1_t_reg[6]), .ZN(
        top_AND_M12_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M12_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_205), .A2(
        top_AND_M12_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M12_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M12_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_169), .A2(top_AND_M12_U1_t_reg[7]), .ZN(
        top_AND_M12_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M12_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M12_U1_OperationInst_q[5]), .A2(
        top_AND_M12_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_232) );
  OR2_X1 top_AND_M12_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M12_U1_OperationInst_q[4]), .A2(
        top_AND_M12_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M12_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M12_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M12_U1_OperationInst_q[7]), .A2(
        top_AND_M12_U1_OperationInst_q[6]), .ZN(
        top_AND_M12_U1_OperationInst_orInst2_n5) );
  OR2_X1 top_XOR_M13_U1_xorInst_U5 ( .A1(top_XOR_M13_U1_xorInst_n12), .A2(
        top_XOR_M13_U1_xorInst_n11), .ZN(top_M13) );
  INV_X1 top_XOR_M13_U1_xorInst_U4 ( .A(top_XOR_M13_U1_xorInst_n10), .ZN(
        top_XOR_M13_U1_xorInst_n11) );
  OR2_X1 top_XOR_M13_U1_xorInst_U3 ( .A1(top_XOR_M13_U1_xorInst_n9), .A2(
        Fresh[7]), .ZN(top_XOR_M13_U1_xorInst_n10) );
  AND2_X1 top_XOR_M13_U1_xorInst_U2 ( .A1(Fresh[7]), .A2(
        top_XOR_M13_U1_xorInst_n9), .ZN(top_XOR_M13_U1_xorInst_n12) );
  INV_X1 top_XOR_M13_U1_xorInst_U1 ( .A(Fresh[6]), .ZN(
        top_XOR_M13_U1_xorInst_n9) );
  AND2_X1 top_XOR_M13_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_229), .A2(
        top_new_AGEMA_signal_232), .ZN(top_XOR_M13_U1_w[0]) );
  AND2_X1 top_XOR_M13_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_230), .A2(
        top_new_AGEMA_signal_231), .ZN(top_XOR_M13_U1_w[1]) );
  AND2_X1 top_XOR_M13_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_230), .A2(
        top_new_AGEMA_signal_232), .ZN(top_XOR_M13_U1_w[2]) );
  AND2_X1 top_XOR_M13_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_229), .A2(
        top_new_AGEMA_signal_231), .ZN(top_XOR_M13_U1_w[3]) );
  OR2_X1 top_XOR_M13_U1_orInst1_U1 ( .A1(top_XOR_M13_U1_w[0]), .A2(
        top_XOR_M13_U1_w[1]), .ZN(top_new_AGEMA_signal_247) );
  OR2_X1 top_XOR_M13_U1_orInst2_U1 ( .A1(top_XOR_M13_U1_w[2]), .A2(
        top_XOR_M13_U1_w[3]), .ZN(top_new_AGEMA_signal_248) );
  INV_X1 top_AND_M14_U1_nonlinearInst_U26 ( .A(top_AND_M14_U1_t[3]), .ZN(
        top_AND_M14_U1_t[7]) );
  OR2_X1 top_AND_M14_U1_nonlinearInst_U25 ( .A1(
        top_AND_M14_U1_nonlinearInst_n64), .A2(
        top_AND_M14_U1_nonlinearInst_n63), .ZN(top_AND_M14_U1_t[3]) );
  INV_X1 top_AND_M14_U1_nonlinearInst_U24 ( .A(
        top_AND_M14_U1_nonlinearInst_n62), .ZN(
        top_AND_M14_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M14_U1_nonlinearInst_U23 ( .A1(
        top_AND_M14_U1_nonlinearInst_n61), .A2(Fresh[8]), .ZN(
        top_AND_M14_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M14_U1_nonlinearInst_U22 ( .A1(Fresh[8]), .A2(
        top_AND_M14_U1_nonlinearInst_n61), .ZN(
        top_AND_M14_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M14_U1_nonlinearInst_U21 ( .A1(top_T2), .A2(top_T10), .ZN(
        top_AND_M14_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M14_U1_nonlinearInst_U20 ( .A(top_AND_M14_U1_t[2]), .ZN(
        top_AND_M14_U1_t[6]) );
  OR2_X1 top_AND_M14_U1_nonlinearInst_U19 ( .A1(
        top_AND_M14_U1_nonlinearInst_n60), .A2(
        top_AND_M14_U1_nonlinearInst_n59), .ZN(top_AND_M14_U1_t[2]) );
  INV_X1 top_AND_M14_U1_nonlinearInst_U18 ( .A(
        top_AND_M14_U1_nonlinearInst_n58), .ZN(
        top_AND_M14_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M14_U1_nonlinearInst_U17 ( .A1(
        top_AND_M14_U1_nonlinearInst_n57), .A2(Fresh[8]), .ZN(
        top_AND_M14_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M14_U1_nonlinearInst_U16 ( .A1(Fresh[8]), .A2(
        top_AND_M14_U1_nonlinearInst_n57), .ZN(
        top_AND_M14_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M14_U1_nonlinearInst_U15 ( .A1(
        top_AND_M14_U1_nonlinearInst_n56), .A2(top_T2), .ZN(
        top_AND_M14_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M14_U1_nonlinearInst_U14 ( .A(top_AND_M14_U1_t[1]), .ZN(
        top_AND_M14_U1_t[5]) );
  OR2_X1 top_AND_M14_U1_nonlinearInst_U13 ( .A1(
        top_AND_M14_U1_nonlinearInst_n55), .A2(
        top_AND_M14_U1_nonlinearInst_n54), .ZN(top_AND_M14_U1_t[1]) );
  AND2_X1 top_AND_M14_U1_nonlinearInst_U12 ( .A1(
        top_AND_M14_U1_nonlinearInst_n53), .A2(
        top_AND_M14_U1_nonlinearInst_n52), .ZN(
        top_AND_M14_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M14_U1_nonlinearInst_U11 ( .A(
        top_AND_M14_U1_nonlinearInst_n51), .ZN(
        top_AND_M14_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M14_U1_nonlinearInst_U10 ( .A1(
        top_AND_M14_U1_nonlinearInst_n52), .A2(
        top_AND_M14_U1_nonlinearInst_n53), .ZN(
        top_AND_M14_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M14_U1_nonlinearInst_U9 ( .A1(top_T2), .A2(
        top_AND_M14_U1_nonlinearInst_n56), .ZN(
        top_AND_M14_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M14_U1_nonlinearInst_U8 ( .A(top_T10), .ZN(
        top_AND_M14_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M14_U1_nonlinearInst_U7 ( .A(top_AND_M14_U1_t[0]), .ZN(
        top_AND_M14_U1_t[4]) );
  OR2_X1 top_AND_M14_U1_nonlinearInst_U6 ( .A1(
        top_AND_M14_U1_nonlinearInst_n50), .A2(
        top_AND_M14_U1_nonlinearInst_n49), .ZN(top_AND_M14_U1_t[0]) );
  AND2_X1 top_AND_M14_U1_nonlinearInst_U5 ( .A1(
        top_AND_M14_U1_nonlinearInst_n48), .A2(
        top_AND_M14_U1_nonlinearInst_n52), .ZN(
        top_AND_M14_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M14_U1_nonlinearInst_U4 ( .A(top_AND_M14_U1_nonlinearInst_n47), .ZN(top_AND_M14_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M14_U1_nonlinearInst_U3 ( .A1(
        top_AND_M14_U1_nonlinearInst_n52), .A2(
        top_AND_M14_U1_nonlinearInst_n48), .ZN(
        top_AND_M14_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M14_U1_nonlinearInst_U2 ( .A1(top_T2), .A2(top_T10), .ZN(
        top_AND_M14_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M14_U1_nonlinearInst_U1 ( .A(Fresh[8]), .ZN(
        top_AND_M14_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M14_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M14_U1_t[0]), .A2(
        top_AND_M14_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M14_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M14_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M14_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M14_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M14_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M14_U1_t_reg[0]) );
  AND2_X1 top_AND_M14_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M14_U1_t[1]), .A2(
        top_AND_M14_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M14_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M14_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M14_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M14_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M14_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M14_U1_t_reg[1]) );
  AND2_X1 top_AND_M14_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M14_U1_t[2]), .A2(
        top_AND_M14_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M14_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M14_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M14_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M14_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M14_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M14_U1_t_reg[2]) );
  AND2_X1 top_AND_M14_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M14_U1_t[3]), .A2(
        top_AND_M14_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M14_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M14_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M14_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M14_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M14_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M14_U1_t_reg[3]) );
  AND2_X1 top_AND_M14_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M14_U1_t[4]), .A2(
        top_AND_M14_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M14_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M14_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M14_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M14_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M14_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M14_U1_t_reg[4]) );
  AND2_X1 top_AND_M14_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M14_U1_t[5]), .A2(
        top_AND_M14_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M14_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M14_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M14_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M14_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M14_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M14_U1_t_reg[5]) );
  AND2_X1 top_AND_M14_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M14_U1_t[6]), .A2(
        top_AND_M14_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M14_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M14_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M14_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M14_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M14_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M14_U1_t_reg[6]) );
  AND2_X1 top_AND_M14_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M14_U1_t[7]), .A2(
        top_AND_M14_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M14_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M14_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M14_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M14_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M14_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M14_U1_t_reg[7]) );
  AND2_X1 top_AND_M14_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_210), .A2(
        top_AND_M14_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M14_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M14_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_164), .A2(top_AND_M14_U1_t_reg[0]), .ZN(
        top_AND_M14_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M14_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_209), .A2(
        top_AND_M14_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M14_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M14_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_164), .A2(top_AND_M14_U1_t_reg[1]), .ZN(
        top_AND_M14_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M14_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_210), .A2(
        top_AND_M14_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M14_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M14_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_163), .A2(top_AND_M14_U1_t_reg[2]), .ZN(
        top_AND_M14_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M14_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_209), .A2(
        top_AND_M14_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M14_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M14_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_163), .A2(top_AND_M14_U1_t_reg[3]), .ZN(
        top_AND_M14_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M14_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M14_U1_OperationInst_q[1]), .A2(
        top_AND_M14_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_249) );
  OR2_X1 top_AND_M14_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M14_U1_OperationInst_q[0]), .A2(
        top_AND_M14_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M14_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M14_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M14_U1_OperationInst_q[3]), .A2(
        top_AND_M14_U1_OperationInst_q[2]), .ZN(
        top_AND_M14_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M14_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_210), .A2(
        top_AND_M14_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M14_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M14_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_164), .A2(top_AND_M14_U1_t_reg[4]), .ZN(
        top_AND_M14_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M14_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_209), .A2(
        top_AND_M14_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M14_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M14_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_164), .A2(top_AND_M14_U1_t_reg[5]), .ZN(
        top_AND_M14_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M14_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_210), .A2(
        top_AND_M14_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M14_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M14_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_163), .A2(top_AND_M14_U1_t_reg[6]), .ZN(
        top_AND_M14_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M14_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_209), .A2(
        top_AND_M14_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M14_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M14_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_163), .A2(top_AND_M14_U1_t_reg[7]), .ZN(
        top_AND_M14_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M14_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M14_U1_OperationInst_q[5]), .A2(
        top_AND_M14_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_250) );
  OR2_X1 top_AND_M14_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M14_U1_OperationInst_q[4]), .A2(
        top_AND_M14_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M14_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M14_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M14_U1_OperationInst_q[7]), .A2(
        top_AND_M14_U1_OperationInst_q[6]), .ZN(
        top_AND_M14_U1_OperationInst_orInst2_n5) );
  OR2_X1 top_XOR_M15_U1_xorInst_U5 ( .A1(top_XOR_M15_U1_xorInst_n12), .A2(
        top_XOR_M15_U1_xorInst_n11), .ZN(top_M15) );
  INV_X1 top_XOR_M15_U1_xorInst_U4 ( .A(top_XOR_M15_U1_xorInst_n10), .ZN(
        top_XOR_M15_U1_xorInst_n11) );
  OR2_X1 top_XOR_M15_U1_xorInst_U3 ( .A1(top_XOR_M15_U1_xorInst_n9), .A2(
        Fresh[8]), .ZN(top_XOR_M15_U1_xorInst_n10) );
  AND2_X1 top_XOR_M15_U1_xorInst_U2 ( .A1(Fresh[8]), .A2(
        top_XOR_M15_U1_xorInst_n9), .ZN(top_XOR_M15_U1_xorInst_n12) );
  INV_X1 top_XOR_M15_U1_xorInst_U1 ( .A(Fresh[6]), .ZN(
        top_XOR_M15_U1_xorInst_n9) );
  AND2_X1 top_XOR_M15_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_229), .A2(
        top_new_AGEMA_signal_250), .ZN(top_XOR_M15_U1_w[0]) );
  AND2_X1 top_XOR_M15_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_230), .A2(
        top_new_AGEMA_signal_249), .ZN(top_XOR_M15_U1_w[1]) );
  AND2_X1 top_XOR_M15_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_230), .A2(
        top_new_AGEMA_signal_250), .ZN(top_XOR_M15_U1_w[2]) );
  AND2_X1 top_XOR_M15_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_229), .A2(
        top_new_AGEMA_signal_249), .ZN(top_XOR_M15_U1_w[3]) );
  OR2_X1 top_XOR_M15_U1_orInst1_U1 ( .A1(top_XOR_M15_U1_w[0]), .A2(
        top_XOR_M15_U1_w[1]), .ZN(top_new_AGEMA_signal_253) );
  OR2_X1 top_XOR_M15_U1_orInst2_U1 ( .A1(top_XOR_M15_U1_w[2]), .A2(
        top_XOR_M15_U1_w[3]), .ZN(top_new_AGEMA_signal_254) );
  OR2_X1 top_XOR_M16_U1_xorInst_U5 ( .A1(top_XOR_M16_U1_xorInst_n12), .A2(
        top_XOR_M16_U1_xorInst_n11), .ZN(top_M16) );
  INV_X1 top_XOR_M16_U1_xorInst_U4 ( .A(top_XOR_M16_U1_xorInst_n10), .ZN(
        top_XOR_M16_U1_xorInst_n11) );
  OR2_X1 top_XOR_M16_U1_xorInst_U3 ( .A1(top_XOR_M16_U1_xorInst_n9), .A2(
        top_M3), .ZN(top_XOR_M16_U1_xorInst_n10) );
  AND2_X1 top_XOR_M16_U1_xorInst_U2 ( .A1(top_M3), .A2(
        top_XOR_M16_U1_xorInst_n9), .ZN(top_XOR_M16_U1_xorInst_n12) );
  INV_X1 top_XOR_M16_U1_xorInst_U1 ( .A(Fresh[1]), .ZN(
        top_XOR_M16_U1_xorInst_n9) );
  AND2_X1 top_XOR_M16_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_237), .A2(
        top_new_AGEMA_signal_240), .ZN(top_XOR_M16_U1_w[0]) );
  AND2_X1 top_XOR_M16_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_238), .A2(
        top_new_AGEMA_signal_239), .ZN(top_XOR_M16_U1_w[1]) );
  AND2_X1 top_XOR_M16_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_238), .A2(
        top_new_AGEMA_signal_240), .ZN(top_XOR_M16_U1_w[2]) );
  AND2_X1 top_XOR_M16_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_237), .A2(
        top_new_AGEMA_signal_239), .ZN(top_XOR_M16_U1_w[3]) );
  OR2_X1 top_XOR_M16_U1_orInst1_U1 ( .A1(top_XOR_M16_U1_w[0]), .A2(
        top_XOR_M16_U1_w[1]), .ZN(top_new_AGEMA_signal_255) );
  OR2_X1 top_XOR_M16_U1_orInst2_U1 ( .A1(top_XOR_M16_U1_w[2]), .A2(
        top_XOR_M16_U1_w[3]), .ZN(top_new_AGEMA_signal_256) );
  OR2_X1 top_XOR_M17_U1_xorInst_U5 ( .A1(top_XOR_M17_U1_xorInst_n12), .A2(
        top_XOR_M17_U1_xorInst_n11), .ZN(top_M17) );
  INV_X1 top_XOR_M17_U1_xorInst_U4 ( .A(top_XOR_M17_U1_xorInst_n10), .ZN(
        top_XOR_M17_U1_xorInst_n11) );
  OR2_X1 top_XOR_M17_U1_xorInst_U3 ( .A1(top_XOR_M17_U1_xorInst_n9), .A2(
        top_M5), .ZN(top_XOR_M17_U1_xorInst_n10) );
  AND2_X1 top_XOR_M17_U1_xorInst_U2 ( .A1(top_M5), .A2(
        top_XOR_M17_U1_xorInst_n9), .ZN(top_XOR_M17_U1_xorInst_n12) );
  INV_X1 top_XOR_M17_U1_xorInst_U1 ( .A(top_T24), .ZN(
        top_XOR_M17_U1_xorInst_n9) );
  AND2_X1 top_XOR_M17_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_233), .A2(
        top_new_AGEMA_signal_242), .ZN(top_XOR_M17_U1_w[0]) );
  AND2_X1 top_XOR_M17_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_234), .A2(
        top_new_AGEMA_signal_241), .ZN(top_XOR_M17_U1_w[1]) );
  AND2_X1 top_XOR_M17_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_234), .A2(
        top_new_AGEMA_signal_242), .ZN(top_XOR_M17_U1_w[2]) );
  AND2_X1 top_XOR_M17_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_233), .A2(
        top_new_AGEMA_signal_241), .ZN(top_XOR_M17_U1_w[3]) );
  OR2_X1 top_XOR_M17_U1_orInst1_U1 ( .A1(top_XOR_M17_U1_w[0]), .A2(
        top_XOR_M17_U1_w[1]), .ZN(top_new_AGEMA_signal_257) );
  OR2_X1 top_XOR_M17_U1_orInst2_U1 ( .A1(top_XOR_M17_U1_w[2]), .A2(
        top_XOR_M17_U1_w[3]), .ZN(top_new_AGEMA_signal_258) );
  OR2_X1 top_XOR_M18_U1_xorInst_U5 ( .A1(top_XOR_M18_U1_xorInst_n12), .A2(
        top_XOR_M18_U1_xorInst_n11), .ZN(top_M18) );
  INV_X1 top_XOR_M18_U1_xorInst_U4 ( .A(top_XOR_M18_U1_xorInst_n10), .ZN(
        top_XOR_M18_U1_xorInst_n11) );
  OR2_X1 top_XOR_M18_U1_xorInst_U3 ( .A1(top_XOR_M18_U1_xorInst_n9), .A2(
        top_M8), .ZN(top_XOR_M18_U1_xorInst_n10) );
  AND2_X1 top_XOR_M18_U1_xorInst_U2 ( .A1(top_M8), .A2(
        top_XOR_M18_U1_xorInst_n9), .ZN(top_XOR_M18_U1_xorInst_n12) );
  INV_X1 top_XOR_M18_U1_xorInst_U1 ( .A(Fresh[4]), .ZN(
        top_XOR_M18_U1_xorInst_n9) );
  AND2_X1 top_XOR_M18_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_227), .A2(
        top_new_AGEMA_signal_244), .ZN(top_XOR_M18_U1_w[0]) );
  AND2_X1 top_XOR_M18_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_228), .A2(
        top_new_AGEMA_signal_243), .ZN(top_XOR_M18_U1_w[1]) );
  AND2_X1 top_XOR_M18_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_228), .A2(
        top_new_AGEMA_signal_244), .ZN(top_XOR_M18_U1_w[2]) );
  AND2_X1 top_XOR_M18_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_227), .A2(
        top_new_AGEMA_signal_243), .ZN(top_XOR_M18_U1_w[3]) );
  OR2_X1 top_XOR_M18_U1_orInst1_U1 ( .A1(top_XOR_M18_U1_w[0]), .A2(
        top_XOR_M18_U1_w[1]), .ZN(top_new_AGEMA_signal_259) );
  OR2_X1 top_XOR_M18_U1_orInst2_U1 ( .A1(top_XOR_M18_U1_w[2]), .A2(
        top_XOR_M18_U1_w[3]), .ZN(top_new_AGEMA_signal_260) );
  OR2_X1 top_XOR_M19_U1_xorInst_U5 ( .A1(top_XOR_M19_U1_xorInst_n12), .A2(
        top_XOR_M19_U1_xorInst_n11), .ZN(top_M19) );
  INV_X1 top_XOR_M19_U1_xorInst_U4 ( .A(top_XOR_M19_U1_xorInst_n10), .ZN(
        top_XOR_M19_U1_xorInst_n11) );
  OR2_X1 top_XOR_M19_U1_xorInst_U3 ( .A1(top_XOR_M19_U1_xorInst_n9), .A2(
        top_M10), .ZN(top_XOR_M19_U1_xorInst_n10) );
  AND2_X1 top_XOR_M19_U1_xorInst_U2 ( .A1(top_M10), .A2(
        top_XOR_M19_U1_xorInst_n9), .ZN(top_XOR_M19_U1_xorInst_n12) );
  INV_X1 top_XOR_M19_U1_xorInst_U1 ( .A(top_M15), .ZN(
        top_XOR_M19_U1_xorInst_n9) );
  AND2_X1 top_XOR_M19_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_253), .A2(
        top_new_AGEMA_signal_252), .ZN(top_XOR_M19_U1_w[0]) );
  AND2_X1 top_XOR_M19_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_254), .A2(
        top_new_AGEMA_signal_251), .ZN(top_XOR_M19_U1_w[1]) );
  AND2_X1 top_XOR_M19_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_254), .A2(
        top_new_AGEMA_signal_252), .ZN(top_XOR_M19_U1_w[2]) );
  AND2_X1 top_XOR_M19_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_253), .A2(
        top_new_AGEMA_signal_251), .ZN(top_XOR_M19_U1_w[3]) );
  OR2_X1 top_XOR_M19_U1_orInst1_U1 ( .A1(top_XOR_M19_U1_w[0]), .A2(
        top_XOR_M19_U1_w[1]), .ZN(top_new_AGEMA_signal_261) );
  OR2_X1 top_XOR_M19_U1_orInst2_U1 ( .A1(top_XOR_M19_U1_w[2]), .A2(
        top_XOR_M19_U1_w[3]), .ZN(top_new_AGEMA_signal_262) );
  OR2_X1 top_XOR_M20_U1_xorInst_U5 ( .A1(top_XOR_M20_U1_xorInst_n12), .A2(
        top_XOR_M20_U1_xorInst_n11), .ZN(top_M20) );
  INV_X1 top_XOR_M20_U1_xorInst_U4 ( .A(top_XOR_M20_U1_xorInst_n10), .ZN(
        top_XOR_M20_U1_xorInst_n11) );
  OR2_X1 top_XOR_M20_U1_xorInst_U3 ( .A1(top_XOR_M20_U1_xorInst_n9), .A2(
        top_M16), .ZN(top_XOR_M20_U1_xorInst_n10) );
  AND2_X1 top_XOR_M20_U1_xorInst_U2 ( .A1(top_M16), .A2(
        top_XOR_M20_U1_xorInst_n9), .ZN(top_XOR_M20_U1_xorInst_n12) );
  INV_X1 top_XOR_M20_U1_xorInst_U1 ( .A(top_M13), .ZN(
        top_XOR_M20_U1_xorInst_n9) );
  AND2_X1 top_XOR_M20_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_247), .A2(
        top_new_AGEMA_signal_256), .ZN(top_XOR_M20_U1_w[0]) );
  AND2_X1 top_XOR_M20_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_248), .A2(
        top_new_AGEMA_signal_255), .ZN(top_XOR_M20_U1_w[1]) );
  AND2_X1 top_XOR_M20_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_248), .A2(
        top_new_AGEMA_signal_256), .ZN(top_XOR_M20_U1_w[2]) );
  AND2_X1 top_XOR_M20_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_247), .A2(
        top_new_AGEMA_signal_255), .ZN(top_XOR_M20_U1_w[3]) );
  OR2_X1 top_XOR_M20_U1_orInst1_U1 ( .A1(top_XOR_M20_U1_w[0]), .A2(
        top_XOR_M20_U1_w[1]), .ZN(top_new_AGEMA_signal_263) );
  OR2_X1 top_XOR_M20_U1_orInst2_U1 ( .A1(top_XOR_M20_U1_w[2]), .A2(
        top_XOR_M20_U1_w[3]), .ZN(top_new_AGEMA_signal_264) );
  OR2_X1 top_XOR_M21_U1_xorInst_U5 ( .A1(top_XOR_M21_U1_xorInst_n12), .A2(
        top_XOR_M21_U1_xorInst_n11), .ZN(top_M21) );
  INV_X1 top_XOR_M21_U1_xorInst_U4 ( .A(top_XOR_M21_U1_xorInst_n10), .ZN(
        top_XOR_M21_U1_xorInst_n11) );
  OR2_X1 top_XOR_M21_U1_xorInst_U3 ( .A1(top_XOR_M21_U1_xorInst_n9), .A2(
        top_M17), .ZN(top_XOR_M21_U1_xorInst_n10) );
  AND2_X1 top_XOR_M21_U1_xorInst_U2 ( .A1(top_M17), .A2(
        top_XOR_M21_U1_xorInst_n9), .ZN(top_XOR_M21_U1_xorInst_n12) );
  INV_X1 top_XOR_M21_U1_xorInst_U1 ( .A(top_M15), .ZN(
        top_XOR_M21_U1_xorInst_n9) );
  AND2_X1 top_XOR_M21_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_253), .A2(
        top_new_AGEMA_signal_258), .ZN(top_XOR_M21_U1_w[0]) );
  AND2_X1 top_XOR_M21_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_254), .A2(
        top_new_AGEMA_signal_257), .ZN(top_XOR_M21_U1_w[1]) );
  AND2_X1 top_XOR_M21_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_254), .A2(
        top_new_AGEMA_signal_258), .ZN(top_XOR_M21_U1_w[2]) );
  AND2_X1 top_XOR_M21_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_253), .A2(
        top_new_AGEMA_signal_257), .ZN(top_XOR_M21_U1_w[3]) );
  OR2_X1 top_XOR_M21_U1_orInst1_U1 ( .A1(top_XOR_M21_U1_w[0]), .A2(
        top_XOR_M21_U1_w[1]), .ZN(top_new_AGEMA_signal_265) );
  OR2_X1 top_XOR_M21_U1_orInst2_U1 ( .A1(top_XOR_M21_U1_w[2]), .A2(
        top_XOR_M21_U1_w[3]), .ZN(top_new_AGEMA_signal_266) );
  OR2_X1 top_XOR_M22_U1_xorInst_U5 ( .A1(top_XOR_M22_U1_xorInst_n12), .A2(
        top_XOR_M22_U1_xorInst_n11), .ZN(top_M22) );
  INV_X1 top_XOR_M22_U1_xorInst_U4 ( .A(top_XOR_M22_U1_xorInst_n10), .ZN(
        top_XOR_M22_U1_xorInst_n11) );
  OR2_X1 top_XOR_M22_U1_xorInst_U3 ( .A1(top_XOR_M22_U1_xorInst_n9), .A2(
        top_M18), .ZN(top_XOR_M22_U1_xorInst_n10) );
  AND2_X1 top_XOR_M22_U1_xorInst_U2 ( .A1(top_M18), .A2(
        top_XOR_M22_U1_xorInst_n9), .ZN(top_XOR_M22_U1_xorInst_n12) );
  INV_X1 top_XOR_M22_U1_xorInst_U1 ( .A(top_M13), .ZN(
        top_XOR_M22_U1_xorInst_n9) );
  AND2_X1 top_XOR_M22_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_247), .A2(
        top_new_AGEMA_signal_260), .ZN(top_XOR_M22_U1_w[0]) );
  AND2_X1 top_XOR_M22_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_248), .A2(
        top_new_AGEMA_signal_259), .ZN(top_XOR_M22_U1_w[1]) );
  AND2_X1 top_XOR_M22_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_248), .A2(
        top_new_AGEMA_signal_260), .ZN(top_XOR_M22_U1_w[2]) );
  AND2_X1 top_XOR_M22_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_247), .A2(
        top_new_AGEMA_signal_259), .ZN(top_XOR_M22_U1_w[3]) );
  OR2_X1 top_XOR_M22_U1_orInst1_U1 ( .A1(top_XOR_M22_U1_w[0]), .A2(
        top_XOR_M22_U1_w[1]), .ZN(top_new_AGEMA_signal_267) );
  OR2_X1 top_XOR_M22_U1_orInst2_U1 ( .A1(top_XOR_M22_U1_w[2]), .A2(
        top_XOR_M22_U1_w[3]), .ZN(top_new_AGEMA_signal_268) );
  OR2_X1 top_XOR_M23_U1_xorInst_U5 ( .A1(top_XOR_M23_U1_xorInst_n12), .A2(
        top_XOR_M23_U1_xorInst_n11), .ZN(top_M23) );
  INV_X1 top_XOR_M23_U1_xorInst_U4 ( .A(top_XOR_M23_U1_xorInst_n10), .ZN(
        top_XOR_M23_U1_xorInst_n11) );
  OR2_X1 top_XOR_M23_U1_xorInst_U3 ( .A1(top_XOR_M23_U1_xorInst_n9), .A2(
        top_M19), .ZN(top_XOR_M23_U1_xorInst_n10) );
  AND2_X1 top_XOR_M23_U1_xorInst_U2 ( .A1(top_M19), .A2(
        top_XOR_M23_U1_xorInst_n9), .ZN(top_XOR_M23_U1_xorInst_n12) );
  INV_X1 top_XOR_M23_U1_xorInst_U1 ( .A(top_T25), .ZN(
        top_XOR_M23_U1_xorInst_n9) );
  AND2_X1 top_XOR_M23_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_235), .A2(
        top_new_AGEMA_signal_262), .ZN(top_XOR_M23_U1_w[0]) );
  AND2_X1 top_XOR_M23_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_236), .A2(
        top_new_AGEMA_signal_261), .ZN(top_XOR_M23_U1_w[1]) );
  AND2_X1 top_XOR_M23_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_236), .A2(
        top_new_AGEMA_signal_262), .ZN(top_XOR_M23_U1_w[2]) );
  AND2_X1 top_XOR_M23_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_235), .A2(
        top_new_AGEMA_signal_261), .ZN(top_XOR_M23_U1_w[3]) );
  OR2_X1 top_XOR_M23_U1_orInst1_U1 ( .A1(top_XOR_M23_U1_w[0]), .A2(
        top_XOR_M23_U1_w[1]), .ZN(top_new_AGEMA_signal_269) );
  OR2_X1 top_XOR_M23_U1_orInst2_U1 ( .A1(top_XOR_M23_U1_w[2]), .A2(
        top_XOR_M23_U1_w[3]), .ZN(top_new_AGEMA_signal_270) );
  OR2_X1 top_XOR_M24_U1_xorInst_U5 ( .A1(top_XOR_M24_U1_xorInst_n12), .A2(
        top_XOR_M24_U1_xorInst_n11), .ZN(top_M24) );
  INV_X1 top_XOR_M24_U1_xorInst_U4 ( .A(top_XOR_M24_U1_xorInst_n10), .ZN(
        top_XOR_M24_U1_xorInst_n11) );
  OR2_X1 top_XOR_M24_U1_xorInst_U3 ( .A1(top_XOR_M24_U1_xorInst_n9), .A2(
        top_M22), .ZN(top_XOR_M24_U1_xorInst_n10) );
  AND2_X1 top_XOR_M24_U1_xorInst_U2 ( .A1(top_M22), .A2(
        top_XOR_M24_U1_xorInst_n9), .ZN(top_XOR_M24_U1_xorInst_n12) );
  INV_X1 top_XOR_M24_U1_xorInst_U1 ( .A(top_M23), .ZN(
        top_XOR_M24_U1_xorInst_n9) );
  AND2_X1 top_XOR_M24_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_269), .A2(
        top_new_AGEMA_signal_268), .ZN(top_XOR_M24_U1_w[0]) );
  AND2_X1 top_XOR_M24_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_270), .A2(
        top_new_AGEMA_signal_267), .ZN(top_XOR_M24_U1_w[1]) );
  AND2_X1 top_XOR_M24_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_270), .A2(
        top_new_AGEMA_signal_268), .ZN(top_XOR_M24_U1_w[2]) );
  AND2_X1 top_XOR_M24_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_269), .A2(
        top_new_AGEMA_signal_267), .ZN(top_XOR_M24_U1_w[3]) );
  OR2_X1 top_XOR_M24_U1_orInst1_U1 ( .A1(top_XOR_M24_U1_w[0]), .A2(
        top_XOR_M24_U1_w[1]), .ZN(top_new_AGEMA_signal_277) );
  OR2_X1 top_XOR_M24_U1_orInst2_U1 ( .A1(top_XOR_M24_U1_w[2]), .A2(
        top_XOR_M24_U1_w[3]), .ZN(top_new_AGEMA_signal_278) );
  INV_X1 top_AND_M25_U1_nonlinearInst_U26 ( .A(top_AND_M25_U1_t[3]), .ZN(
        top_AND_M25_U1_t[7]) );
  OR2_X1 top_AND_M25_U1_nonlinearInst_U25 ( .A1(
        top_AND_M25_U1_nonlinearInst_n64), .A2(
        top_AND_M25_U1_nonlinearInst_n63), .ZN(top_AND_M25_U1_t[3]) );
  INV_X1 top_AND_M25_U1_nonlinearInst_U24 ( .A(
        top_AND_M25_U1_nonlinearInst_n62), .ZN(
        top_AND_M25_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M25_U1_nonlinearInst_U23 ( .A1(
        top_AND_M25_U1_nonlinearInst_n61), .A2(Fresh[9]), .ZN(
        top_AND_M25_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M25_U1_nonlinearInst_U22 ( .A1(Fresh[9]), .A2(
        top_AND_M25_U1_nonlinearInst_n61), .ZN(
        top_AND_M25_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M25_U1_nonlinearInst_U21 ( .A1(top_M22), .A2(top_M20), .ZN(
        top_AND_M25_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M25_U1_nonlinearInst_U20 ( .A(top_AND_M25_U1_t[2]), .ZN(
        top_AND_M25_U1_t[6]) );
  OR2_X1 top_AND_M25_U1_nonlinearInst_U19 ( .A1(
        top_AND_M25_U1_nonlinearInst_n60), .A2(
        top_AND_M25_U1_nonlinearInst_n59), .ZN(top_AND_M25_U1_t[2]) );
  INV_X1 top_AND_M25_U1_nonlinearInst_U18 ( .A(
        top_AND_M25_U1_nonlinearInst_n58), .ZN(
        top_AND_M25_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M25_U1_nonlinearInst_U17 ( .A1(
        top_AND_M25_U1_nonlinearInst_n57), .A2(Fresh[9]), .ZN(
        top_AND_M25_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M25_U1_nonlinearInst_U16 ( .A1(Fresh[9]), .A2(
        top_AND_M25_U1_nonlinearInst_n57), .ZN(
        top_AND_M25_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M25_U1_nonlinearInst_U15 ( .A1(
        top_AND_M25_U1_nonlinearInst_n56), .A2(top_M22), .ZN(
        top_AND_M25_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M25_U1_nonlinearInst_U14 ( .A(top_AND_M25_U1_t[1]), .ZN(
        top_AND_M25_U1_t[5]) );
  OR2_X1 top_AND_M25_U1_nonlinearInst_U13 ( .A1(
        top_AND_M25_U1_nonlinearInst_n55), .A2(
        top_AND_M25_U1_nonlinearInst_n54), .ZN(top_AND_M25_U1_t[1]) );
  AND2_X1 top_AND_M25_U1_nonlinearInst_U12 ( .A1(
        top_AND_M25_U1_nonlinearInst_n53), .A2(
        top_AND_M25_U1_nonlinearInst_n52), .ZN(
        top_AND_M25_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M25_U1_nonlinearInst_U11 ( .A(
        top_AND_M25_U1_nonlinearInst_n51), .ZN(
        top_AND_M25_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M25_U1_nonlinearInst_U10 ( .A1(
        top_AND_M25_U1_nonlinearInst_n52), .A2(
        top_AND_M25_U1_nonlinearInst_n53), .ZN(
        top_AND_M25_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M25_U1_nonlinearInst_U9 ( .A1(top_M22), .A2(
        top_AND_M25_U1_nonlinearInst_n56), .ZN(
        top_AND_M25_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M25_U1_nonlinearInst_U8 ( .A(top_M20), .ZN(
        top_AND_M25_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M25_U1_nonlinearInst_U7 ( .A(top_AND_M25_U1_t[0]), .ZN(
        top_AND_M25_U1_t[4]) );
  OR2_X1 top_AND_M25_U1_nonlinearInst_U6 ( .A1(
        top_AND_M25_U1_nonlinearInst_n50), .A2(
        top_AND_M25_U1_nonlinearInst_n49), .ZN(top_AND_M25_U1_t[0]) );
  AND2_X1 top_AND_M25_U1_nonlinearInst_U5 ( .A1(
        top_AND_M25_U1_nonlinearInst_n48), .A2(
        top_AND_M25_U1_nonlinearInst_n52), .ZN(
        top_AND_M25_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M25_U1_nonlinearInst_U4 ( .A(top_AND_M25_U1_nonlinearInst_n47), .ZN(top_AND_M25_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M25_U1_nonlinearInst_U3 ( .A1(
        top_AND_M25_U1_nonlinearInst_n52), .A2(
        top_AND_M25_U1_nonlinearInst_n48), .ZN(
        top_AND_M25_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M25_U1_nonlinearInst_U2 ( .A1(top_M22), .A2(top_M20), .ZN(
        top_AND_M25_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M25_U1_nonlinearInst_U1 ( .A(Fresh[9]), .ZN(
        top_AND_M25_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M25_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M25_U1_t[0]), .A2(
        top_AND_M25_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M25_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M25_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M25_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M25_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M25_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M25_U1_t_reg[0]) );
  AND2_X1 top_AND_M25_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M25_U1_t[1]), .A2(
        top_AND_M25_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M25_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M25_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M25_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M25_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M25_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M25_U1_t_reg[1]) );
  AND2_X1 top_AND_M25_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M25_U1_t[2]), .A2(
        top_AND_M25_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M25_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M25_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M25_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M25_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M25_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M25_U1_t_reg[2]) );
  AND2_X1 top_AND_M25_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M25_U1_t[3]), .A2(
        top_AND_M25_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M25_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M25_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M25_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M25_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M25_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M25_U1_t_reg[3]) );
  AND2_X1 top_AND_M25_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M25_U1_t[4]), .A2(
        top_AND_M25_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M25_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M25_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M25_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M25_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M25_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M25_U1_t_reg[4]) );
  AND2_X1 top_AND_M25_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M25_U1_t[5]), .A2(
        top_AND_M25_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M25_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M25_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M25_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M25_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M25_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M25_U1_t_reg[5]) );
  AND2_X1 top_AND_M25_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M25_U1_t[6]), .A2(
        top_AND_M25_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M25_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M25_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M25_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M25_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M25_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M25_U1_t_reg[6]) );
  AND2_X1 top_AND_M25_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M25_U1_t[7]), .A2(
        top_AND_M25_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M25_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M25_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M25_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M25_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M25_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M25_U1_t_reg[7]) );
  AND2_X1 top_AND_M25_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_264), .A2(
        top_AND_M25_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M25_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M25_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_268), .A2(top_AND_M25_U1_t_reg[0]), .ZN(
        top_AND_M25_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M25_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_263), .A2(
        top_AND_M25_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M25_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M25_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_268), .A2(top_AND_M25_U1_t_reg[1]), .ZN(
        top_AND_M25_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M25_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_264), .A2(
        top_AND_M25_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M25_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M25_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_267), .A2(top_AND_M25_U1_t_reg[2]), .ZN(
        top_AND_M25_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M25_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_263), .A2(
        top_AND_M25_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M25_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M25_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_267), .A2(top_AND_M25_U1_t_reg[3]), .ZN(
        top_AND_M25_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M25_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M25_U1_OperationInst_q[1]), .A2(
        top_AND_M25_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_271) );
  OR2_X1 top_AND_M25_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M25_U1_OperationInst_q[0]), .A2(
        top_AND_M25_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M25_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M25_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M25_U1_OperationInst_q[3]), .A2(
        top_AND_M25_U1_OperationInst_q[2]), .ZN(
        top_AND_M25_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M25_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_264), .A2(
        top_AND_M25_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M25_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M25_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_268), .A2(top_AND_M25_U1_t_reg[4]), .ZN(
        top_AND_M25_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M25_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_263), .A2(
        top_AND_M25_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M25_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M25_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_268), .A2(top_AND_M25_U1_t_reg[5]), .ZN(
        top_AND_M25_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M25_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_264), .A2(
        top_AND_M25_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M25_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M25_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_267), .A2(top_AND_M25_U1_t_reg[6]), .ZN(
        top_AND_M25_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M25_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_263), .A2(
        top_AND_M25_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M25_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M25_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_267), .A2(top_AND_M25_U1_t_reg[7]), .ZN(
        top_AND_M25_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M25_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M25_U1_OperationInst_q[5]), .A2(
        top_AND_M25_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_272) );
  OR2_X1 top_AND_M25_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M25_U1_OperationInst_q[4]), .A2(
        top_AND_M25_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M25_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M25_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M25_U1_OperationInst_q[7]), .A2(
        top_AND_M25_U1_OperationInst_q[6]), .ZN(
        top_AND_M25_U1_OperationInst_orInst2_n5) );
  OR2_X1 top_XOR_M26_U1_xorInst_U5 ( .A1(top_XOR_M26_U1_xorInst_n12), .A2(
        top_XOR_M26_U1_xorInst_n11), .ZN(top_M26) );
  INV_X1 top_XOR_M26_U1_xorInst_U4 ( .A(top_XOR_M26_U1_xorInst_n10), .ZN(
        top_XOR_M26_U1_xorInst_n11) );
  OR2_X1 top_XOR_M26_U1_xorInst_U3 ( .A1(top_XOR_M26_U1_xorInst_n9), .A2(
        top_M21), .ZN(top_XOR_M26_U1_xorInst_n10) );
  AND2_X1 top_XOR_M26_U1_xorInst_U2 ( .A1(top_M21), .A2(
        top_XOR_M26_U1_xorInst_n9), .ZN(top_XOR_M26_U1_xorInst_n12) );
  INV_X1 top_XOR_M26_U1_xorInst_U1 ( .A(Fresh[9]), .ZN(
        top_XOR_M26_U1_xorInst_n9) );
  AND2_X1 top_XOR_M26_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_271), .A2(
        top_new_AGEMA_signal_266), .ZN(top_XOR_M26_U1_w[0]) );
  AND2_X1 top_XOR_M26_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_272), .A2(
        top_new_AGEMA_signal_265), .ZN(top_XOR_M26_U1_w[1]) );
  AND2_X1 top_XOR_M26_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_272), .A2(
        top_new_AGEMA_signal_266), .ZN(top_XOR_M26_U1_w[2]) );
  AND2_X1 top_XOR_M26_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_271), .A2(
        top_new_AGEMA_signal_265), .ZN(top_XOR_M26_U1_w[3]) );
  OR2_X1 top_XOR_M26_U1_orInst1_U1 ( .A1(top_XOR_M26_U1_w[0]), .A2(
        top_XOR_M26_U1_w[1]), .ZN(top_new_AGEMA_signal_279) );
  OR2_X1 top_XOR_M26_U1_orInst2_U1 ( .A1(top_XOR_M26_U1_w[2]), .A2(
        top_XOR_M26_U1_w[3]), .ZN(top_new_AGEMA_signal_280) );
  OR2_X1 top_XOR_M27_U1_xorInst_U5 ( .A1(top_XOR_M27_U1_xorInst_n12), .A2(
        top_XOR_M27_U1_xorInst_n11), .ZN(top_M27) );
  INV_X1 top_XOR_M27_U1_xorInst_U4 ( .A(top_XOR_M27_U1_xorInst_n10), .ZN(
        top_XOR_M27_U1_xorInst_n11) );
  OR2_X1 top_XOR_M27_U1_xorInst_U3 ( .A1(top_XOR_M27_U1_xorInst_n9), .A2(
        top_M20), .ZN(top_XOR_M27_U1_xorInst_n10) );
  AND2_X1 top_XOR_M27_U1_xorInst_U2 ( .A1(top_M20), .A2(
        top_XOR_M27_U1_xorInst_n9), .ZN(top_XOR_M27_U1_xorInst_n12) );
  INV_X1 top_XOR_M27_U1_xorInst_U1 ( .A(top_M21), .ZN(
        top_XOR_M27_U1_xorInst_n9) );
  AND2_X1 top_XOR_M27_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_265), .A2(
        top_new_AGEMA_signal_264), .ZN(top_XOR_M27_U1_w[0]) );
  AND2_X1 top_XOR_M27_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_266), .A2(
        top_new_AGEMA_signal_263), .ZN(top_XOR_M27_U1_w[1]) );
  AND2_X1 top_XOR_M27_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_266), .A2(
        top_new_AGEMA_signal_264), .ZN(top_XOR_M27_U1_w[2]) );
  AND2_X1 top_XOR_M27_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_265), .A2(
        top_new_AGEMA_signal_263), .ZN(top_XOR_M27_U1_w[3]) );
  OR2_X1 top_XOR_M27_U1_orInst1_U1 ( .A1(top_XOR_M27_U1_w[0]), .A2(
        top_XOR_M27_U1_w[1]), .ZN(top_new_AGEMA_signal_273) );
  OR2_X1 top_XOR_M27_U1_orInst2_U1 ( .A1(top_XOR_M27_U1_w[2]), .A2(
        top_XOR_M27_U1_w[3]), .ZN(top_new_AGEMA_signal_274) );
  OR2_X1 top_XOR_M28_U1_xorInst_U5 ( .A1(top_XOR_M28_U1_xorInst_n12), .A2(
        top_XOR_M28_U1_xorInst_n11), .ZN(top_M28) );
  INV_X1 top_XOR_M28_U1_xorInst_U4 ( .A(top_XOR_M28_U1_xorInst_n10), .ZN(
        top_XOR_M28_U1_xorInst_n11) );
  OR2_X1 top_XOR_M28_U1_xorInst_U3 ( .A1(top_XOR_M28_U1_xorInst_n9), .A2(
        top_M23), .ZN(top_XOR_M28_U1_xorInst_n10) );
  AND2_X1 top_XOR_M28_U1_xorInst_U2 ( .A1(top_M23), .A2(
        top_XOR_M28_U1_xorInst_n9), .ZN(top_XOR_M28_U1_xorInst_n12) );
  INV_X1 top_XOR_M28_U1_xorInst_U1 ( .A(Fresh[9]), .ZN(
        top_XOR_M28_U1_xorInst_n9) );
  AND2_X1 top_XOR_M28_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_271), .A2(
        top_new_AGEMA_signal_270), .ZN(top_XOR_M28_U1_w[0]) );
  AND2_X1 top_XOR_M28_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_272), .A2(
        top_new_AGEMA_signal_269), .ZN(top_XOR_M28_U1_w[1]) );
  AND2_X1 top_XOR_M28_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_272), .A2(
        top_new_AGEMA_signal_270), .ZN(top_XOR_M28_U1_w[2]) );
  AND2_X1 top_XOR_M28_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_271), .A2(
        top_new_AGEMA_signal_269), .ZN(top_XOR_M28_U1_w[3]) );
  OR2_X1 top_XOR_M28_U1_orInst1_U1 ( .A1(top_XOR_M28_U1_w[0]), .A2(
        top_XOR_M28_U1_w[1]), .ZN(top_new_AGEMA_signal_281) );
  OR2_X1 top_XOR_M28_U1_orInst2_U1 ( .A1(top_XOR_M28_U1_w[2]), .A2(
        top_XOR_M28_U1_w[3]), .ZN(top_new_AGEMA_signal_282) );
  INV_X1 top_AND_M29_U1_nonlinearInst_U26 ( .A(top_AND_M29_U1_t[3]), .ZN(
        top_AND_M29_U1_t[7]) );
  OR2_X1 top_AND_M29_U1_nonlinearInst_U25 ( .A1(
        top_AND_M29_U1_nonlinearInst_n64), .A2(
        top_AND_M29_U1_nonlinearInst_n63), .ZN(top_AND_M29_U1_t[3]) );
  INV_X1 top_AND_M29_U1_nonlinearInst_U24 ( .A(
        top_AND_M29_U1_nonlinearInst_n62), .ZN(
        top_AND_M29_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M29_U1_nonlinearInst_U23 ( .A1(
        top_AND_M29_U1_nonlinearInst_n61), .A2(Fresh[10]), .ZN(
        top_AND_M29_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M29_U1_nonlinearInst_U22 ( .A1(Fresh[10]), .A2(
        top_AND_M29_U1_nonlinearInst_n61), .ZN(
        top_AND_M29_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M29_U1_nonlinearInst_U21 ( .A1(top_M28), .A2(top_M27), .ZN(
        top_AND_M29_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M29_U1_nonlinearInst_U20 ( .A(top_AND_M29_U1_t[2]), .ZN(
        top_AND_M29_U1_t[6]) );
  OR2_X1 top_AND_M29_U1_nonlinearInst_U19 ( .A1(
        top_AND_M29_U1_nonlinearInst_n60), .A2(
        top_AND_M29_U1_nonlinearInst_n59), .ZN(top_AND_M29_U1_t[2]) );
  INV_X1 top_AND_M29_U1_nonlinearInst_U18 ( .A(
        top_AND_M29_U1_nonlinearInst_n58), .ZN(
        top_AND_M29_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M29_U1_nonlinearInst_U17 ( .A1(
        top_AND_M29_U1_nonlinearInst_n57), .A2(Fresh[10]), .ZN(
        top_AND_M29_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M29_U1_nonlinearInst_U16 ( .A1(Fresh[10]), .A2(
        top_AND_M29_U1_nonlinearInst_n57), .ZN(
        top_AND_M29_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M29_U1_nonlinearInst_U15 ( .A1(
        top_AND_M29_U1_nonlinearInst_n56), .A2(top_M28), .ZN(
        top_AND_M29_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M29_U1_nonlinearInst_U14 ( .A(top_AND_M29_U1_t[1]), .ZN(
        top_AND_M29_U1_t[5]) );
  OR2_X1 top_AND_M29_U1_nonlinearInst_U13 ( .A1(
        top_AND_M29_U1_nonlinearInst_n55), .A2(
        top_AND_M29_U1_nonlinearInst_n54), .ZN(top_AND_M29_U1_t[1]) );
  AND2_X1 top_AND_M29_U1_nonlinearInst_U12 ( .A1(
        top_AND_M29_U1_nonlinearInst_n53), .A2(
        top_AND_M29_U1_nonlinearInst_n52), .ZN(
        top_AND_M29_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M29_U1_nonlinearInst_U11 ( .A(
        top_AND_M29_U1_nonlinearInst_n51), .ZN(
        top_AND_M29_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M29_U1_nonlinearInst_U10 ( .A1(
        top_AND_M29_U1_nonlinearInst_n52), .A2(
        top_AND_M29_U1_nonlinearInst_n53), .ZN(
        top_AND_M29_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M29_U1_nonlinearInst_U9 ( .A1(top_M28), .A2(
        top_AND_M29_U1_nonlinearInst_n56), .ZN(
        top_AND_M29_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M29_U1_nonlinearInst_U8 ( .A(top_M27), .ZN(
        top_AND_M29_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M29_U1_nonlinearInst_U7 ( .A(top_AND_M29_U1_t[0]), .ZN(
        top_AND_M29_U1_t[4]) );
  OR2_X1 top_AND_M29_U1_nonlinearInst_U6 ( .A1(
        top_AND_M29_U1_nonlinearInst_n50), .A2(
        top_AND_M29_U1_nonlinearInst_n49), .ZN(top_AND_M29_U1_t[0]) );
  AND2_X1 top_AND_M29_U1_nonlinearInst_U5 ( .A1(
        top_AND_M29_U1_nonlinearInst_n48), .A2(
        top_AND_M29_U1_nonlinearInst_n52), .ZN(
        top_AND_M29_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M29_U1_nonlinearInst_U4 ( .A(top_AND_M29_U1_nonlinearInst_n47), .ZN(top_AND_M29_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M29_U1_nonlinearInst_U3 ( .A1(
        top_AND_M29_U1_nonlinearInst_n52), .A2(
        top_AND_M29_U1_nonlinearInst_n48), .ZN(
        top_AND_M29_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M29_U1_nonlinearInst_U2 ( .A1(top_M28), .A2(top_M27), .ZN(
        top_AND_M29_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M29_U1_nonlinearInst_U1 ( .A(Fresh[10]), .ZN(
        top_AND_M29_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M29_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M29_U1_t[0]), .A2(
        top_AND_M29_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M29_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M29_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M29_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M29_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M29_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M29_U1_t_reg[0]) );
  AND2_X1 top_AND_M29_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M29_U1_t[1]), .A2(
        top_AND_M29_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M29_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M29_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M29_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M29_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M29_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M29_U1_t_reg[1]) );
  AND2_X1 top_AND_M29_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M29_U1_t[2]), .A2(
        top_AND_M29_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M29_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M29_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M29_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M29_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M29_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M29_U1_t_reg[2]) );
  AND2_X1 top_AND_M29_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M29_U1_t[3]), .A2(
        top_AND_M29_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M29_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M29_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M29_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M29_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M29_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M29_U1_t_reg[3]) );
  AND2_X1 top_AND_M29_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M29_U1_t[4]), .A2(
        top_AND_M29_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M29_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M29_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M29_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M29_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M29_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M29_U1_t_reg[4]) );
  AND2_X1 top_AND_M29_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M29_U1_t[5]), .A2(
        top_AND_M29_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M29_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M29_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M29_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M29_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M29_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M29_U1_t_reg[5]) );
  AND2_X1 top_AND_M29_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M29_U1_t[6]), .A2(
        top_AND_M29_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M29_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M29_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M29_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M29_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M29_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M29_U1_t_reg[6]) );
  AND2_X1 top_AND_M29_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M29_U1_t[7]), .A2(
        top_AND_M29_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M29_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M29_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M29_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M29_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M29_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M29_U1_t_reg[7]) );
  AND2_X1 top_AND_M29_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_274), .A2(
        top_AND_M29_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M29_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M29_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_282), .A2(top_AND_M29_U1_t_reg[0]), .ZN(
        top_AND_M29_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M29_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_273), .A2(
        top_AND_M29_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M29_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M29_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_282), .A2(top_AND_M29_U1_t_reg[1]), .ZN(
        top_AND_M29_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M29_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_274), .A2(
        top_AND_M29_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M29_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M29_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_281), .A2(top_AND_M29_U1_t_reg[2]), .ZN(
        top_AND_M29_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M29_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_273), .A2(
        top_AND_M29_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M29_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M29_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_281), .A2(top_AND_M29_U1_t_reg[3]), .ZN(
        top_AND_M29_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M29_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M29_U1_OperationInst_q[1]), .A2(
        top_AND_M29_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_287) );
  OR2_X1 top_AND_M29_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M29_U1_OperationInst_q[0]), .A2(
        top_AND_M29_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M29_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M29_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M29_U1_OperationInst_q[3]), .A2(
        top_AND_M29_U1_OperationInst_q[2]), .ZN(
        top_AND_M29_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M29_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_274), .A2(
        top_AND_M29_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M29_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M29_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_282), .A2(top_AND_M29_U1_t_reg[4]), .ZN(
        top_AND_M29_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M29_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_273), .A2(
        top_AND_M29_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M29_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M29_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_282), .A2(top_AND_M29_U1_t_reg[5]), .ZN(
        top_AND_M29_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M29_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_274), .A2(
        top_AND_M29_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M29_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M29_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_281), .A2(top_AND_M29_U1_t_reg[6]), .ZN(
        top_AND_M29_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M29_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_273), .A2(
        top_AND_M29_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M29_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M29_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_281), .A2(top_AND_M29_U1_t_reg[7]), .ZN(
        top_AND_M29_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M29_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M29_U1_OperationInst_q[5]), .A2(
        top_AND_M29_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_288) );
  OR2_X1 top_AND_M29_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M29_U1_OperationInst_q[4]), .A2(
        top_AND_M29_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M29_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M29_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M29_U1_OperationInst_q[7]), .A2(
        top_AND_M29_U1_OperationInst_q[6]), .ZN(
        top_AND_M29_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M30_U1_nonlinearInst_U26 ( .A(top_AND_M30_U1_t[3]), .ZN(
        top_AND_M30_U1_t[7]) );
  OR2_X1 top_AND_M30_U1_nonlinearInst_U25 ( .A1(
        top_AND_M30_U1_nonlinearInst_n64), .A2(
        top_AND_M30_U1_nonlinearInst_n63), .ZN(top_AND_M30_U1_t[3]) );
  INV_X1 top_AND_M30_U1_nonlinearInst_U24 ( .A(
        top_AND_M30_U1_nonlinearInst_n62), .ZN(
        top_AND_M30_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M30_U1_nonlinearInst_U23 ( .A1(
        top_AND_M30_U1_nonlinearInst_n61), .A2(Fresh[11]), .ZN(
        top_AND_M30_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M30_U1_nonlinearInst_U22 ( .A1(Fresh[11]), .A2(
        top_AND_M30_U1_nonlinearInst_n61), .ZN(
        top_AND_M30_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M30_U1_nonlinearInst_U21 ( .A1(top_M26), .A2(top_M24), .ZN(
        top_AND_M30_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M30_U1_nonlinearInst_U20 ( .A(top_AND_M30_U1_t[2]), .ZN(
        top_AND_M30_U1_t[6]) );
  OR2_X1 top_AND_M30_U1_nonlinearInst_U19 ( .A1(
        top_AND_M30_U1_nonlinearInst_n60), .A2(
        top_AND_M30_U1_nonlinearInst_n59), .ZN(top_AND_M30_U1_t[2]) );
  INV_X1 top_AND_M30_U1_nonlinearInst_U18 ( .A(
        top_AND_M30_U1_nonlinearInst_n58), .ZN(
        top_AND_M30_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M30_U1_nonlinearInst_U17 ( .A1(
        top_AND_M30_U1_nonlinearInst_n57), .A2(Fresh[11]), .ZN(
        top_AND_M30_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M30_U1_nonlinearInst_U16 ( .A1(Fresh[11]), .A2(
        top_AND_M30_U1_nonlinearInst_n57), .ZN(
        top_AND_M30_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M30_U1_nonlinearInst_U15 ( .A1(
        top_AND_M30_U1_nonlinearInst_n56), .A2(top_M26), .ZN(
        top_AND_M30_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M30_U1_nonlinearInst_U14 ( .A(top_AND_M30_U1_t[1]), .ZN(
        top_AND_M30_U1_t[5]) );
  OR2_X1 top_AND_M30_U1_nonlinearInst_U13 ( .A1(
        top_AND_M30_U1_nonlinearInst_n55), .A2(
        top_AND_M30_U1_nonlinearInst_n54), .ZN(top_AND_M30_U1_t[1]) );
  AND2_X1 top_AND_M30_U1_nonlinearInst_U12 ( .A1(
        top_AND_M30_U1_nonlinearInst_n53), .A2(
        top_AND_M30_U1_nonlinearInst_n52), .ZN(
        top_AND_M30_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M30_U1_nonlinearInst_U11 ( .A(
        top_AND_M30_U1_nonlinearInst_n51), .ZN(
        top_AND_M30_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M30_U1_nonlinearInst_U10 ( .A1(
        top_AND_M30_U1_nonlinearInst_n52), .A2(
        top_AND_M30_U1_nonlinearInst_n53), .ZN(
        top_AND_M30_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M30_U1_nonlinearInst_U9 ( .A1(top_M26), .A2(
        top_AND_M30_U1_nonlinearInst_n56), .ZN(
        top_AND_M30_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M30_U1_nonlinearInst_U8 ( .A(top_M24), .ZN(
        top_AND_M30_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M30_U1_nonlinearInst_U7 ( .A(top_AND_M30_U1_t[0]), .ZN(
        top_AND_M30_U1_t[4]) );
  OR2_X1 top_AND_M30_U1_nonlinearInst_U6 ( .A1(
        top_AND_M30_U1_nonlinearInst_n50), .A2(
        top_AND_M30_U1_nonlinearInst_n49), .ZN(top_AND_M30_U1_t[0]) );
  AND2_X1 top_AND_M30_U1_nonlinearInst_U5 ( .A1(
        top_AND_M30_U1_nonlinearInst_n48), .A2(
        top_AND_M30_U1_nonlinearInst_n52), .ZN(
        top_AND_M30_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M30_U1_nonlinearInst_U4 ( .A(top_AND_M30_U1_nonlinearInst_n47), .ZN(top_AND_M30_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M30_U1_nonlinearInst_U3 ( .A1(
        top_AND_M30_U1_nonlinearInst_n52), .A2(
        top_AND_M30_U1_nonlinearInst_n48), .ZN(
        top_AND_M30_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M30_U1_nonlinearInst_U2 ( .A1(top_M26), .A2(top_M24), .ZN(
        top_AND_M30_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M30_U1_nonlinearInst_U1 ( .A(Fresh[11]), .ZN(
        top_AND_M30_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M30_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M30_U1_t[0]), .A2(
        top_AND_M30_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M30_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M30_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M30_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M30_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M30_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M30_U1_t_reg[0]) );
  AND2_X1 top_AND_M30_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M30_U1_t[1]), .A2(
        top_AND_M30_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M30_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M30_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M30_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M30_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M30_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M30_U1_t_reg[1]) );
  AND2_X1 top_AND_M30_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M30_U1_t[2]), .A2(
        top_AND_M30_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M30_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M30_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M30_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M30_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M30_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M30_U1_t_reg[2]) );
  AND2_X1 top_AND_M30_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M30_U1_t[3]), .A2(
        top_AND_M30_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M30_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M30_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M30_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M30_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M30_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M30_U1_t_reg[3]) );
  AND2_X1 top_AND_M30_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M30_U1_t[4]), .A2(
        top_AND_M30_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M30_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M30_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M30_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M30_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M30_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M30_U1_t_reg[4]) );
  AND2_X1 top_AND_M30_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M30_U1_t[5]), .A2(
        top_AND_M30_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M30_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M30_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M30_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M30_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M30_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M30_U1_t_reg[5]) );
  AND2_X1 top_AND_M30_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M30_U1_t[6]), .A2(
        top_AND_M30_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M30_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M30_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M30_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M30_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M30_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M30_U1_t_reg[6]) );
  AND2_X1 top_AND_M30_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M30_U1_t[7]), .A2(
        top_AND_M30_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M30_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M30_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M30_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M30_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M30_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M30_U1_t_reg[7]) );
  AND2_X1 top_AND_M30_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_278), .A2(
        top_AND_M30_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M30_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M30_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_280), .A2(top_AND_M30_U1_t_reg[0]), .ZN(
        top_AND_M30_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M30_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_277), .A2(
        top_AND_M30_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M30_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M30_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_280), .A2(top_AND_M30_U1_t_reg[1]), .ZN(
        top_AND_M30_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M30_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_278), .A2(
        top_AND_M30_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M30_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M30_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_279), .A2(top_AND_M30_U1_t_reg[2]), .ZN(
        top_AND_M30_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M30_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_277), .A2(
        top_AND_M30_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M30_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M30_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_279), .A2(top_AND_M30_U1_t_reg[3]), .ZN(
        top_AND_M30_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M30_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M30_U1_OperationInst_q[1]), .A2(
        top_AND_M30_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_289) );
  OR2_X1 top_AND_M30_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M30_U1_OperationInst_q[0]), .A2(
        top_AND_M30_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M30_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M30_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M30_U1_OperationInst_q[3]), .A2(
        top_AND_M30_U1_OperationInst_q[2]), .ZN(
        top_AND_M30_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M30_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_278), .A2(
        top_AND_M30_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M30_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M30_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_280), .A2(top_AND_M30_U1_t_reg[4]), .ZN(
        top_AND_M30_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M30_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_277), .A2(
        top_AND_M30_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M30_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M30_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_280), .A2(top_AND_M30_U1_t_reg[5]), .ZN(
        top_AND_M30_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M30_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_278), .A2(
        top_AND_M30_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M30_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M30_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_279), .A2(top_AND_M30_U1_t_reg[6]), .ZN(
        top_AND_M30_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M30_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_277), .A2(
        top_AND_M30_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M30_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M30_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_279), .A2(top_AND_M30_U1_t_reg[7]), .ZN(
        top_AND_M30_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M30_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M30_U1_OperationInst_q[5]), .A2(
        top_AND_M30_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_290) );
  OR2_X1 top_AND_M30_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M30_U1_OperationInst_q[4]), .A2(
        top_AND_M30_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M30_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M30_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M30_U1_OperationInst_q[7]), .A2(
        top_AND_M30_U1_OperationInst_q[6]), .ZN(
        top_AND_M30_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M31_U1_nonlinearInst_U26 ( .A(top_AND_M31_U1_t[3]), .ZN(
        top_AND_M31_U1_t[7]) );
  OR2_X1 top_AND_M31_U1_nonlinearInst_U25 ( .A1(
        top_AND_M31_U1_nonlinearInst_n64), .A2(
        top_AND_M31_U1_nonlinearInst_n63), .ZN(top_AND_M31_U1_t[3]) );
  INV_X1 top_AND_M31_U1_nonlinearInst_U24 ( .A(
        top_AND_M31_U1_nonlinearInst_n62), .ZN(
        top_AND_M31_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M31_U1_nonlinearInst_U23 ( .A1(
        top_AND_M31_U1_nonlinearInst_n61), .A2(Fresh[12]), .ZN(
        top_AND_M31_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M31_U1_nonlinearInst_U22 ( .A1(Fresh[12]), .A2(
        top_AND_M31_U1_nonlinearInst_n61), .ZN(
        top_AND_M31_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M31_U1_nonlinearInst_U21 ( .A1(top_M20), .A2(top_M23), .ZN(
        top_AND_M31_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M31_U1_nonlinearInst_U20 ( .A(top_AND_M31_U1_t[2]), .ZN(
        top_AND_M31_U1_t[6]) );
  OR2_X1 top_AND_M31_U1_nonlinearInst_U19 ( .A1(
        top_AND_M31_U1_nonlinearInst_n60), .A2(
        top_AND_M31_U1_nonlinearInst_n59), .ZN(top_AND_M31_U1_t[2]) );
  INV_X1 top_AND_M31_U1_nonlinearInst_U18 ( .A(
        top_AND_M31_U1_nonlinearInst_n58), .ZN(
        top_AND_M31_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M31_U1_nonlinearInst_U17 ( .A1(
        top_AND_M31_U1_nonlinearInst_n57), .A2(Fresh[12]), .ZN(
        top_AND_M31_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M31_U1_nonlinearInst_U16 ( .A1(Fresh[12]), .A2(
        top_AND_M31_U1_nonlinearInst_n57), .ZN(
        top_AND_M31_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M31_U1_nonlinearInst_U15 ( .A1(
        top_AND_M31_U1_nonlinearInst_n56), .A2(top_M20), .ZN(
        top_AND_M31_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M31_U1_nonlinearInst_U14 ( .A(top_AND_M31_U1_t[1]), .ZN(
        top_AND_M31_U1_t[5]) );
  OR2_X1 top_AND_M31_U1_nonlinearInst_U13 ( .A1(
        top_AND_M31_U1_nonlinearInst_n55), .A2(
        top_AND_M31_U1_nonlinearInst_n54), .ZN(top_AND_M31_U1_t[1]) );
  AND2_X1 top_AND_M31_U1_nonlinearInst_U12 ( .A1(
        top_AND_M31_U1_nonlinearInst_n53), .A2(
        top_AND_M31_U1_nonlinearInst_n52), .ZN(
        top_AND_M31_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M31_U1_nonlinearInst_U11 ( .A(
        top_AND_M31_U1_nonlinearInst_n51), .ZN(
        top_AND_M31_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M31_U1_nonlinearInst_U10 ( .A1(
        top_AND_M31_U1_nonlinearInst_n52), .A2(
        top_AND_M31_U1_nonlinearInst_n53), .ZN(
        top_AND_M31_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M31_U1_nonlinearInst_U9 ( .A1(top_M20), .A2(
        top_AND_M31_U1_nonlinearInst_n56), .ZN(
        top_AND_M31_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M31_U1_nonlinearInst_U8 ( .A(top_M23), .ZN(
        top_AND_M31_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M31_U1_nonlinearInst_U7 ( .A(top_AND_M31_U1_t[0]), .ZN(
        top_AND_M31_U1_t[4]) );
  OR2_X1 top_AND_M31_U1_nonlinearInst_U6 ( .A1(
        top_AND_M31_U1_nonlinearInst_n50), .A2(
        top_AND_M31_U1_nonlinearInst_n49), .ZN(top_AND_M31_U1_t[0]) );
  AND2_X1 top_AND_M31_U1_nonlinearInst_U5 ( .A1(
        top_AND_M31_U1_nonlinearInst_n48), .A2(
        top_AND_M31_U1_nonlinearInst_n52), .ZN(
        top_AND_M31_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M31_U1_nonlinearInst_U4 ( .A(top_AND_M31_U1_nonlinearInst_n47), .ZN(top_AND_M31_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M31_U1_nonlinearInst_U3 ( .A1(
        top_AND_M31_U1_nonlinearInst_n52), .A2(
        top_AND_M31_U1_nonlinearInst_n48), .ZN(
        top_AND_M31_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M31_U1_nonlinearInst_U2 ( .A1(top_M20), .A2(top_M23), .ZN(
        top_AND_M31_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M31_U1_nonlinearInst_U1 ( .A(Fresh[12]), .ZN(
        top_AND_M31_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M31_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M31_U1_t[0]), .A2(
        top_AND_M31_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M31_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M31_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M31_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M31_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M31_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M31_U1_t_reg[0]) );
  AND2_X1 top_AND_M31_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M31_U1_t[1]), .A2(
        top_AND_M31_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M31_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M31_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M31_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M31_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M31_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M31_U1_t_reg[1]) );
  AND2_X1 top_AND_M31_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M31_U1_t[2]), .A2(
        top_AND_M31_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M31_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M31_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M31_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M31_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M31_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M31_U1_t_reg[2]) );
  AND2_X1 top_AND_M31_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M31_U1_t[3]), .A2(
        top_AND_M31_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M31_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M31_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M31_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M31_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M31_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M31_U1_t_reg[3]) );
  AND2_X1 top_AND_M31_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M31_U1_t[4]), .A2(
        top_AND_M31_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M31_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M31_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M31_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M31_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M31_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M31_U1_t_reg[4]) );
  AND2_X1 top_AND_M31_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M31_U1_t[5]), .A2(
        top_AND_M31_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M31_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M31_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M31_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M31_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M31_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M31_U1_t_reg[5]) );
  AND2_X1 top_AND_M31_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M31_U1_t[6]), .A2(
        top_AND_M31_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M31_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M31_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M31_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M31_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M31_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M31_U1_t_reg[6]) );
  AND2_X1 top_AND_M31_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M31_U1_t[7]), .A2(
        top_AND_M31_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M31_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M31_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M31_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M31_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M31_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M31_U1_t_reg[7]) );
  AND2_X1 top_AND_M31_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_270), .A2(
        top_AND_M31_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M31_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M31_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_264), .A2(top_AND_M31_U1_t_reg[0]), .ZN(
        top_AND_M31_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M31_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_269), .A2(
        top_AND_M31_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M31_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M31_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_264), .A2(top_AND_M31_U1_t_reg[1]), .ZN(
        top_AND_M31_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M31_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_270), .A2(
        top_AND_M31_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M31_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M31_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_263), .A2(top_AND_M31_U1_t_reg[2]), .ZN(
        top_AND_M31_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M31_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_269), .A2(
        top_AND_M31_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M31_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M31_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_263), .A2(top_AND_M31_U1_t_reg[3]), .ZN(
        top_AND_M31_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M31_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M31_U1_OperationInst_q[1]), .A2(
        top_AND_M31_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_283) );
  OR2_X1 top_AND_M31_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M31_U1_OperationInst_q[0]), .A2(
        top_AND_M31_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M31_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M31_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M31_U1_OperationInst_q[3]), .A2(
        top_AND_M31_U1_OperationInst_q[2]), .ZN(
        top_AND_M31_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M31_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_270), .A2(
        top_AND_M31_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M31_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M31_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_264), .A2(top_AND_M31_U1_t_reg[4]), .ZN(
        top_AND_M31_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M31_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_269), .A2(
        top_AND_M31_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M31_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M31_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_264), .A2(top_AND_M31_U1_t_reg[5]), .ZN(
        top_AND_M31_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M31_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_270), .A2(
        top_AND_M31_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M31_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M31_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_263), .A2(top_AND_M31_U1_t_reg[6]), .ZN(
        top_AND_M31_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M31_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_269), .A2(
        top_AND_M31_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M31_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M31_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_263), .A2(top_AND_M31_U1_t_reg[7]), .ZN(
        top_AND_M31_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M31_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M31_U1_OperationInst_q[5]), .A2(
        top_AND_M31_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_284) );
  OR2_X1 top_AND_M31_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M31_U1_OperationInst_q[4]), .A2(
        top_AND_M31_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M31_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M31_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M31_U1_OperationInst_q[7]), .A2(
        top_AND_M31_U1_OperationInst_q[6]), .ZN(
        top_AND_M31_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M32_U1_nonlinearInst_U26 ( .A(top_AND_M32_U1_t[3]), .ZN(
        top_AND_M32_U1_t[7]) );
  OR2_X1 top_AND_M32_U1_nonlinearInst_U25 ( .A1(
        top_AND_M32_U1_nonlinearInst_n64), .A2(
        top_AND_M32_U1_nonlinearInst_n63), .ZN(top_AND_M32_U1_t[3]) );
  INV_X1 top_AND_M32_U1_nonlinearInst_U24 ( .A(
        top_AND_M32_U1_nonlinearInst_n62), .ZN(
        top_AND_M32_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M32_U1_nonlinearInst_U23 ( .A1(
        top_AND_M32_U1_nonlinearInst_n61), .A2(Fresh[13]), .ZN(
        top_AND_M32_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M32_U1_nonlinearInst_U22 ( .A1(Fresh[13]), .A2(
        top_AND_M32_U1_nonlinearInst_n61), .ZN(
        top_AND_M32_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M32_U1_nonlinearInst_U21 ( .A1(top_M27), .A2(Fresh[12]), .ZN(
        top_AND_M32_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M32_U1_nonlinearInst_U20 ( .A(top_AND_M32_U1_t[2]), .ZN(
        top_AND_M32_U1_t[6]) );
  OR2_X1 top_AND_M32_U1_nonlinearInst_U19 ( .A1(
        top_AND_M32_U1_nonlinearInst_n60), .A2(
        top_AND_M32_U1_nonlinearInst_n59), .ZN(top_AND_M32_U1_t[2]) );
  INV_X1 top_AND_M32_U1_nonlinearInst_U18 ( .A(
        top_AND_M32_U1_nonlinearInst_n58), .ZN(
        top_AND_M32_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M32_U1_nonlinearInst_U17 ( .A1(
        top_AND_M32_U1_nonlinearInst_n57), .A2(Fresh[13]), .ZN(
        top_AND_M32_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M32_U1_nonlinearInst_U16 ( .A1(Fresh[13]), .A2(
        top_AND_M32_U1_nonlinearInst_n57), .ZN(
        top_AND_M32_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M32_U1_nonlinearInst_U15 ( .A1(
        top_AND_M32_U1_nonlinearInst_n56), .A2(top_M27), .ZN(
        top_AND_M32_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M32_U1_nonlinearInst_U14 ( .A(top_AND_M32_U1_t[1]), .ZN(
        top_AND_M32_U1_t[5]) );
  OR2_X1 top_AND_M32_U1_nonlinearInst_U13 ( .A1(
        top_AND_M32_U1_nonlinearInst_n55), .A2(
        top_AND_M32_U1_nonlinearInst_n54), .ZN(top_AND_M32_U1_t[1]) );
  AND2_X1 top_AND_M32_U1_nonlinearInst_U12 ( .A1(
        top_AND_M32_U1_nonlinearInst_n53), .A2(
        top_AND_M32_U1_nonlinearInst_n52), .ZN(
        top_AND_M32_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M32_U1_nonlinearInst_U11 ( .A(
        top_AND_M32_U1_nonlinearInst_n51), .ZN(
        top_AND_M32_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M32_U1_nonlinearInst_U10 ( .A1(
        top_AND_M32_U1_nonlinearInst_n52), .A2(
        top_AND_M32_U1_nonlinearInst_n53), .ZN(
        top_AND_M32_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M32_U1_nonlinearInst_U9 ( .A1(top_M27), .A2(
        top_AND_M32_U1_nonlinearInst_n56), .ZN(
        top_AND_M32_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M32_U1_nonlinearInst_U8 ( .A(Fresh[12]), .ZN(
        top_AND_M32_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M32_U1_nonlinearInst_U7 ( .A(top_AND_M32_U1_t[0]), .ZN(
        top_AND_M32_U1_t[4]) );
  OR2_X1 top_AND_M32_U1_nonlinearInst_U6 ( .A1(
        top_AND_M32_U1_nonlinearInst_n50), .A2(
        top_AND_M32_U1_nonlinearInst_n49), .ZN(top_AND_M32_U1_t[0]) );
  AND2_X1 top_AND_M32_U1_nonlinearInst_U5 ( .A1(
        top_AND_M32_U1_nonlinearInst_n48), .A2(
        top_AND_M32_U1_nonlinearInst_n52), .ZN(
        top_AND_M32_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M32_U1_nonlinearInst_U4 ( .A(top_AND_M32_U1_nonlinearInst_n47), .ZN(top_AND_M32_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M32_U1_nonlinearInst_U3 ( .A1(
        top_AND_M32_U1_nonlinearInst_n52), .A2(
        top_AND_M32_U1_nonlinearInst_n48), .ZN(
        top_AND_M32_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M32_U1_nonlinearInst_U2 ( .A1(top_M27), .A2(Fresh[12]), .ZN(
        top_AND_M32_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M32_U1_nonlinearInst_U1 ( .A(Fresh[13]), .ZN(
        top_AND_M32_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M32_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M32_U1_t[0]), .A2(
        top_AND_M32_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M32_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M32_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M32_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M32_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M32_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M32_U1_t_reg[0]) );
  AND2_X1 top_AND_M32_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M32_U1_t[1]), .A2(
        top_AND_M32_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M32_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M32_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M32_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M32_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M32_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M32_U1_t_reg[1]) );
  AND2_X1 top_AND_M32_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M32_U1_t[2]), .A2(
        top_AND_M32_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M32_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M32_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M32_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M32_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M32_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M32_U1_t_reg[2]) );
  AND2_X1 top_AND_M32_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M32_U1_t[3]), .A2(
        top_AND_M32_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M32_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M32_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M32_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M32_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M32_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M32_U1_t_reg[3]) );
  AND2_X1 top_AND_M32_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M32_U1_t[4]), .A2(
        top_AND_M32_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M32_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M32_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M32_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M32_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M32_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M32_U1_t_reg[4]) );
  AND2_X1 top_AND_M32_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M32_U1_t[5]), .A2(
        top_AND_M32_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M32_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M32_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M32_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M32_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M32_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M32_U1_t_reg[5]) );
  AND2_X1 top_AND_M32_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M32_U1_t[6]), .A2(
        top_AND_M32_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M32_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M32_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M32_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M32_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M32_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M32_U1_t_reg[6]) );
  AND2_X1 top_AND_M32_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M32_U1_t[7]), .A2(
        top_AND_M32_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M32_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M32_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M32_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M32_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M32_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M32_U1_t_reg[7]) );
  AND2_X1 top_AND_M32_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_284), .A2(
        top_AND_M32_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M32_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M32_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_274), .A2(top_AND_M32_U1_t_reg[0]), .ZN(
        top_AND_M32_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M32_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_283), .A2(
        top_AND_M32_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M32_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M32_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_274), .A2(top_AND_M32_U1_t_reg[1]), .ZN(
        top_AND_M32_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M32_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_284), .A2(
        top_AND_M32_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M32_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M32_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_273), .A2(top_AND_M32_U1_t_reg[2]), .ZN(
        top_AND_M32_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M32_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_283), .A2(
        top_AND_M32_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M32_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M32_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_273), .A2(top_AND_M32_U1_t_reg[3]), .ZN(
        top_AND_M32_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M32_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M32_U1_OperationInst_q[1]), .A2(
        top_AND_M32_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_291) );
  OR2_X1 top_AND_M32_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M32_U1_OperationInst_q[0]), .A2(
        top_AND_M32_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M32_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M32_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M32_U1_OperationInst_q[3]), .A2(
        top_AND_M32_U1_OperationInst_q[2]), .ZN(
        top_AND_M32_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M32_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_284), .A2(
        top_AND_M32_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M32_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M32_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_274), .A2(top_AND_M32_U1_t_reg[4]), .ZN(
        top_AND_M32_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M32_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_283), .A2(
        top_AND_M32_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M32_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M32_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_274), .A2(top_AND_M32_U1_t_reg[5]), .ZN(
        top_AND_M32_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M32_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_284), .A2(
        top_AND_M32_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M32_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M32_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_273), .A2(top_AND_M32_U1_t_reg[6]), .ZN(
        top_AND_M32_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M32_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_283), .A2(
        top_AND_M32_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M32_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M32_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_273), .A2(top_AND_M32_U1_t_reg[7]), .ZN(
        top_AND_M32_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M32_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M32_U1_OperationInst_q[5]), .A2(
        top_AND_M32_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_292) );
  OR2_X1 top_AND_M32_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M32_U1_OperationInst_q[4]), .A2(
        top_AND_M32_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M32_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M32_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M32_U1_OperationInst_q[7]), .A2(
        top_AND_M32_U1_OperationInst_q[6]), .ZN(
        top_AND_M32_U1_OperationInst_orInst2_n5) );
  OR2_X1 top_XOR_M33_U1_xorInst_U5 ( .A1(top_XOR_M33_U1_xorInst_n12), .A2(
        top_XOR_M33_U1_xorInst_n11), .ZN(top_M33) );
  INV_X1 top_XOR_M33_U1_xorInst_U4 ( .A(top_XOR_M33_U1_xorInst_n10), .ZN(
        top_XOR_M33_U1_xorInst_n11) );
  OR2_X1 top_XOR_M33_U1_xorInst_U3 ( .A1(top_XOR_M33_U1_xorInst_n9), .A2(
        top_M27), .ZN(top_XOR_M33_U1_xorInst_n10) );
  AND2_X1 top_XOR_M33_U1_xorInst_U2 ( .A1(top_M27), .A2(
        top_XOR_M33_U1_xorInst_n9), .ZN(top_XOR_M33_U1_xorInst_n12) );
  INV_X1 top_XOR_M33_U1_xorInst_U1 ( .A(Fresh[9]), .ZN(
        top_XOR_M33_U1_xorInst_n9) );
  AND2_X1 top_XOR_M33_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_271), .A2(
        top_new_AGEMA_signal_274), .ZN(top_XOR_M33_U1_w[0]) );
  AND2_X1 top_XOR_M33_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_272), .A2(
        top_new_AGEMA_signal_273), .ZN(top_XOR_M33_U1_w[1]) );
  AND2_X1 top_XOR_M33_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_272), .A2(
        top_new_AGEMA_signal_274), .ZN(top_XOR_M33_U1_w[2]) );
  AND2_X1 top_XOR_M33_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_271), .A2(
        top_new_AGEMA_signal_273), .ZN(top_XOR_M33_U1_w[3]) );
  OR2_X1 top_XOR_M33_U1_orInst1_U1 ( .A1(top_XOR_M33_U1_w[0]), .A2(
        top_XOR_M33_U1_w[1]), .ZN(top_new_AGEMA_signal_285) );
  OR2_X1 top_XOR_M33_U1_orInst2_U1 ( .A1(top_XOR_M33_U1_w[2]), .A2(
        top_XOR_M33_U1_w[3]), .ZN(top_new_AGEMA_signal_286) );
  INV_X1 top_AND_M34_U1_nonlinearInst_U26 ( .A(top_AND_M34_U1_t[3]), .ZN(
        top_AND_M34_U1_t[7]) );
  OR2_X1 top_AND_M34_U1_nonlinearInst_U25 ( .A1(
        top_AND_M34_U1_nonlinearInst_n64), .A2(
        top_AND_M34_U1_nonlinearInst_n63), .ZN(top_AND_M34_U1_t[3]) );
  INV_X1 top_AND_M34_U1_nonlinearInst_U24 ( .A(
        top_AND_M34_U1_nonlinearInst_n62), .ZN(
        top_AND_M34_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M34_U1_nonlinearInst_U23 ( .A1(
        top_AND_M34_U1_nonlinearInst_n61), .A2(Fresh[14]), .ZN(
        top_AND_M34_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M34_U1_nonlinearInst_U22 ( .A1(Fresh[14]), .A2(
        top_AND_M34_U1_nonlinearInst_n61), .ZN(
        top_AND_M34_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M34_U1_nonlinearInst_U21 ( .A1(top_M21), .A2(top_M22), .ZN(
        top_AND_M34_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M34_U1_nonlinearInst_U20 ( .A(top_AND_M34_U1_t[2]), .ZN(
        top_AND_M34_U1_t[6]) );
  OR2_X1 top_AND_M34_U1_nonlinearInst_U19 ( .A1(
        top_AND_M34_U1_nonlinearInst_n60), .A2(
        top_AND_M34_U1_nonlinearInst_n59), .ZN(top_AND_M34_U1_t[2]) );
  INV_X1 top_AND_M34_U1_nonlinearInst_U18 ( .A(
        top_AND_M34_U1_nonlinearInst_n58), .ZN(
        top_AND_M34_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M34_U1_nonlinearInst_U17 ( .A1(
        top_AND_M34_U1_nonlinearInst_n57), .A2(Fresh[14]), .ZN(
        top_AND_M34_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M34_U1_nonlinearInst_U16 ( .A1(Fresh[14]), .A2(
        top_AND_M34_U1_nonlinearInst_n57), .ZN(
        top_AND_M34_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M34_U1_nonlinearInst_U15 ( .A1(
        top_AND_M34_U1_nonlinearInst_n56), .A2(top_M21), .ZN(
        top_AND_M34_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M34_U1_nonlinearInst_U14 ( .A(top_AND_M34_U1_t[1]), .ZN(
        top_AND_M34_U1_t[5]) );
  OR2_X1 top_AND_M34_U1_nonlinearInst_U13 ( .A1(
        top_AND_M34_U1_nonlinearInst_n55), .A2(
        top_AND_M34_U1_nonlinearInst_n54), .ZN(top_AND_M34_U1_t[1]) );
  AND2_X1 top_AND_M34_U1_nonlinearInst_U12 ( .A1(
        top_AND_M34_U1_nonlinearInst_n53), .A2(
        top_AND_M34_U1_nonlinearInst_n52), .ZN(
        top_AND_M34_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M34_U1_nonlinearInst_U11 ( .A(
        top_AND_M34_U1_nonlinearInst_n51), .ZN(
        top_AND_M34_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M34_U1_nonlinearInst_U10 ( .A1(
        top_AND_M34_U1_nonlinearInst_n52), .A2(
        top_AND_M34_U1_nonlinearInst_n53), .ZN(
        top_AND_M34_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M34_U1_nonlinearInst_U9 ( .A1(top_M21), .A2(
        top_AND_M34_U1_nonlinearInst_n56), .ZN(
        top_AND_M34_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M34_U1_nonlinearInst_U8 ( .A(top_M22), .ZN(
        top_AND_M34_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M34_U1_nonlinearInst_U7 ( .A(top_AND_M34_U1_t[0]), .ZN(
        top_AND_M34_U1_t[4]) );
  OR2_X1 top_AND_M34_U1_nonlinearInst_U6 ( .A1(
        top_AND_M34_U1_nonlinearInst_n50), .A2(
        top_AND_M34_U1_nonlinearInst_n49), .ZN(top_AND_M34_U1_t[0]) );
  AND2_X1 top_AND_M34_U1_nonlinearInst_U5 ( .A1(
        top_AND_M34_U1_nonlinearInst_n48), .A2(
        top_AND_M34_U1_nonlinearInst_n52), .ZN(
        top_AND_M34_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M34_U1_nonlinearInst_U4 ( .A(top_AND_M34_U1_nonlinearInst_n47), .ZN(top_AND_M34_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M34_U1_nonlinearInst_U3 ( .A1(
        top_AND_M34_U1_nonlinearInst_n52), .A2(
        top_AND_M34_U1_nonlinearInst_n48), .ZN(
        top_AND_M34_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M34_U1_nonlinearInst_U2 ( .A1(top_M21), .A2(top_M22), .ZN(
        top_AND_M34_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M34_U1_nonlinearInst_U1 ( .A(Fresh[14]), .ZN(
        top_AND_M34_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M34_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M34_U1_t[0]), .A2(
        top_AND_M34_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M34_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M34_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M34_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M34_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M34_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M34_U1_t_reg[0]) );
  AND2_X1 top_AND_M34_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M34_U1_t[1]), .A2(
        top_AND_M34_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M34_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M34_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M34_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M34_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M34_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M34_U1_t_reg[1]) );
  AND2_X1 top_AND_M34_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M34_U1_t[2]), .A2(
        top_AND_M34_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M34_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M34_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M34_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M34_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M34_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M34_U1_t_reg[2]) );
  AND2_X1 top_AND_M34_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M34_U1_t[3]), .A2(
        top_AND_M34_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M34_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M34_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M34_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M34_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M34_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M34_U1_t_reg[3]) );
  AND2_X1 top_AND_M34_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M34_U1_t[4]), .A2(
        top_AND_M34_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M34_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M34_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M34_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M34_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M34_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M34_U1_t_reg[4]) );
  AND2_X1 top_AND_M34_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M34_U1_t[5]), .A2(
        top_AND_M34_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M34_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M34_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M34_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M34_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M34_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M34_U1_t_reg[5]) );
  AND2_X1 top_AND_M34_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M34_U1_t[6]), .A2(
        top_AND_M34_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M34_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M34_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M34_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M34_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M34_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M34_U1_t_reg[6]) );
  AND2_X1 top_AND_M34_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M34_U1_t[7]), .A2(
        top_AND_M34_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M34_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M34_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M34_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M34_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M34_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M34_U1_t_reg[7]) );
  AND2_X1 top_AND_M34_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_268), .A2(
        top_AND_M34_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M34_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M34_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_266), .A2(top_AND_M34_U1_t_reg[0]), .ZN(
        top_AND_M34_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M34_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_267), .A2(
        top_AND_M34_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M34_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M34_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_266), .A2(top_AND_M34_U1_t_reg[1]), .ZN(
        top_AND_M34_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M34_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_268), .A2(
        top_AND_M34_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M34_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M34_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_265), .A2(top_AND_M34_U1_t_reg[2]), .ZN(
        top_AND_M34_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M34_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_267), .A2(
        top_AND_M34_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M34_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M34_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_265), .A2(top_AND_M34_U1_t_reg[3]), .ZN(
        top_AND_M34_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M34_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M34_U1_OperationInst_q[1]), .A2(
        top_AND_M34_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_275) );
  OR2_X1 top_AND_M34_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M34_U1_OperationInst_q[0]), .A2(
        top_AND_M34_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M34_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M34_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M34_U1_OperationInst_q[3]), .A2(
        top_AND_M34_U1_OperationInst_q[2]), .ZN(
        top_AND_M34_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M34_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_268), .A2(
        top_AND_M34_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M34_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M34_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_266), .A2(top_AND_M34_U1_t_reg[4]), .ZN(
        top_AND_M34_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M34_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_267), .A2(
        top_AND_M34_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M34_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M34_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_266), .A2(top_AND_M34_U1_t_reg[5]), .ZN(
        top_AND_M34_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M34_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_268), .A2(
        top_AND_M34_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M34_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M34_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_265), .A2(top_AND_M34_U1_t_reg[6]), .ZN(
        top_AND_M34_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M34_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_267), .A2(
        top_AND_M34_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M34_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M34_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_265), .A2(top_AND_M34_U1_t_reg[7]), .ZN(
        top_AND_M34_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M34_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M34_U1_OperationInst_q[5]), .A2(
        top_AND_M34_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_276) );
  OR2_X1 top_AND_M34_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M34_U1_OperationInst_q[4]), .A2(
        top_AND_M34_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M34_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M34_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M34_U1_OperationInst_q[7]), .A2(
        top_AND_M34_U1_OperationInst_q[6]), .ZN(
        top_AND_M34_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M35_U1_nonlinearInst_U26 ( .A(top_AND_M35_U1_t[3]), .ZN(
        top_AND_M35_U1_t[7]) );
  OR2_X1 top_AND_M35_U1_nonlinearInst_U25 ( .A1(
        top_AND_M35_U1_nonlinearInst_n64), .A2(
        top_AND_M35_U1_nonlinearInst_n63), .ZN(top_AND_M35_U1_t[3]) );
  INV_X1 top_AND_M35_U1_nonlinearInst_U24 ( .A(
        top_AND_M35_U1_nonlinearInst_n62), .ZN(
        top_AND_M35_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M35_U1_nonlinearInst_U23 ( .A1(
        top_AND_M35_U1_nonlinearInst_n61), .A2(Fresh[15]), .ZN(
        top_AND_M35_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M35_U1_nonlinearInst_U22 ( .A1(Fresh[15]), .A2(
        top_AND_M35_U1_nonlinearInst_n61), .ZN(
        top_AND_M35_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M35_U1_nonlinearInst_U21 ( .A1(top_M24), .A2(Fresh[14]), .ZN(
        top_AND_M35_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M35_U1_nonlinearInst_U20 ( .A(top_AND_M35_U1_t[1]), .ZN(
        top_AND_M35_U1_t[5]) );
  OR2_X1 top_AND_M35_U1_nonlinearInst_U19 ( .A1(
        top_AND_M35_U1_nonlinearInst_n60), .A2(
        top_AND_M35_U1_nonlinearInst_n59), .ZN(top_AND_M35_U1_t[1]) );
  AND2_X1 top_AND_M35_U1_nonlinearInst_U18 ( .A1(
        top_AND_M35_U1_nonlinearInst_n58), .A2(
        top_AND_M35_U1_nonlinearInst_n57), .ZN(
        top_AND_M35_U1_nonlinearInst_n59) );
  INV_X1 top_AND_M35_U1_nonlinearInst_U17 ( .A(
        top_AND_M35_U1_nonlinearInst_n56), .ZN(
        top_AND_M35_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M35_U1_nonlinearInst_U16 ( .A1(
        top_AND_M35_U1_nonlinearInst_n57), .A2(
        top_AND_M35_U1_nonlinearInst_n58), .ZN(
        top_AND_M35_U1_nonlinearInst_n56) );
  AND2_X1 top_AND_M35_U1_nonlinearInst_U15 ( .A1(top_M24), .A2(
        top_AND_M35_U1_nonlinearInst_n55), .ZN(
        top_AND_M35_U1_nonlinearInst_n58) );
  INV_X1 top_AND_M35_U1_nonlinearInst_U14 ( .A(top_AND_M35_U1_t[0]), .ZN(
        top_AND_M35_U1_t[4]) );
  OR2_X1 top_AND_M35_U1_nonlinearInst_U13 ( .A1(
        top_AND_M35_U1_nonlinearInst_n54), .A2(
        top_AND_M35_U1_nonlinearInst_n53), .ZN(top_AND_M35_U1_t[0]) );
  AND2_X1 top_AND_M35_U1_nonlinearInst_U12 ( .A1(
        top_AND_M35_U1_nonlinearInst_n52), .A2(
        top_AND_M35_U1_nonlinearInst_n57), .ZN(
        top_AND_M35_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M35_U1_nonlinearInst_U11 ( .A(
        top_AND_M35_U1_nonlinearInst_n51), .ZN(
        top_AND_M35_U1_nonlinearInst_n54) );
  OR2_X1 top_AND_M35_U1_nonlinearInst_U10 ( .A1(
        top_AND_M35_U1_nonlinearInst_n57), .A2(
        top_AND_M35_U1_nonlinearInst_n52), .ZN(
        top_AND_M35_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M35_U1_nonlinearInst_U9 ( .A1(top_M24), .A2(Fresh[14]), .ZN(
        top_AND_M35_U1_nonlinearInst_n52) );
  INV_X1 top_AND_M35_U1_nonlinearInst_U8 ( .A(Fresh[15]), .ZN(
        top_AND_M35_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M35_U1_nonlinearInst_U7 ( .A(top_AND_M35_U1_t[2]), .ZN(
        top_AND_M35_U1_t[6]) );
  OR2_X1 top_AND_M35_U1_nonlinearInst_U6 ( .A1(
        top_AND_M35_U1_nonlinearInst_n50), .A2(
        top_AND_M35_U1_nonlinearInst_n49), .ZN(top_AND_M35_U1_t[2]) );
  INV_X1 top_AND_M35_U1_nonlinearInst_U5 ( .A(top_AND_M35_U1_nonlinearInst_n48), .ZN(top_AND_M35_U1_nonlinearInst_n49) );
  OR2_X1 top_AND_M35_U1_nonlinearInst_U4 ( .A1(
        top_AND_M35_U1_nonlinearInst_n47), .A2(Fresh[15]), .ZN(
        top_AND_M35_U1_nonlinearInst_n48) );
  AND2_X1 top_AND_M35_U1_nonlinearInst_U3 ( .A1(Fresh[15]), .A2(
        top_AND_M35_U1_nonlinearInst_n47), .ZN(
        top_AND_M35_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M35_U1_nonlinearInst_U2 ( .A1(
        top_AND_M35_U1_nonlinearInst_n55), .A2(top_M24), .ZN(
        top_AND_M35_U1_nonlinearInst_n47) );
  INV_X1 top_AND_M35_U1_nonlinearInst_U1 ( .A(Fresh[14]), .ZN(
        top_AND_M35_U1_nonlinearInst_n55) );
  AND2_X1 top_AND_M35_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M35_U1_t[0]), .A2(
        top_AND_M35_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M35_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M35_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M35_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M35_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M35_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M35_U1_t_reg[0]) );
  AND2_X1 top_AND_M35_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M35_U1_t[1]), .A2(
        top_AND_M35_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M35_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M35_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M35_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M35_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M35_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M35_U1_t_reg[1]) );
  AND2_X1 top_AND_M35_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M35_U1_t[2]), .A2(
        top_AND_M35_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M35_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M35_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M35_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M35_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M35_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M35_U1_t_reg[2]) );
  AND2_X1 top_AND_M35_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M35_U1_t[3]), .A2(
        top_AND_M35_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M35_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M35_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M35_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M35_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M35_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M35_U1_t_reg[3]) );
  AND2_X1 top_AND_M35_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M35_U1_t[4]), .A2(
        top_AND_M35_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M35_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M35_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M35_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M35_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M35_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M35_U1_t_reg[4]) );
  AND2_X1 top_AND_M35_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M35_U1_t[5]), .A2(
        top_AND_M35_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M35_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M35_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M35_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M35_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M35_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M35_U1_t_reg[5]) );
  AND2_X1 top_AND_M35_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M35_U1_t[6]), .A2(
        top_AND_M35_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M35_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M35_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M35_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M35_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M35_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M35_U1_t_reg[6]) );
  AND2_X1 top_AND_M35_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M35_U1_t[7]), .A2(
        top_AND_M35_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M35_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M35_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M35_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M35_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M35_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M35_U1_t_reg[7]) );
  AND2_X1 top_AND_M35_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_276), .A2(
        top_AND_M35_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M35_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M35_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_278), .A2(top_AND_M35_U1_t_reg[0]), .ZN(
        top_AND_M35_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M35_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_275), .A2(
        top_AND_M35_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M35_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M35_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_278), .A2(top_AND_M35_U1_t_reg[1]), .ZN(
        top_AND_M35_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M35_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_276), .A2(
        top_AND_M35_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M35_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M35_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_277), .A2(top_AND_M35_U1_t_reg[2]), .ZN(
        top_AND_M35_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M35_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_275), .A2(
        top_AND_M35_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M35_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M35_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_277), .A2(top_AND_M35_U1_t_reg[3]), .ZN(
        top_AND_M35_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M35_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M35_U1_OperationInst_q[1]), .A2(
        top_AND_M35_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_293) );
  OR2_X1 top_AND_M35_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M35_U1_OperationInst_q[0]), .A2(
        top_AND_M35_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M35_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M35_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M35_U1_OperationInst_q[3]), .A2(
        top_AND_M35_U1_OperationInst_q[2]), .ZN(
        top_AND_M35_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M35_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_276), .A2(
        top_AND_M35_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M35_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M35_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_278), .A2(top_AND_M35_U1_t_reg[4]), .ZN(
        top_AND_M35_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M35_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_275), .A2(
        top_AND_M35_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M35_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M35_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_278), .A2(top_AND_M35_U1_t_reg[5]), .ZN(
        top_AND_M35_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M35_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_276), .A2(
        top_AND_M35_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M35_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M35_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_277), .A2(top_AND_M35_U1_t_reg[6]), .ZN(
        top_AND_M35_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M35_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_275), .A2(
        top_AND_M35_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M35_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M35_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_277), .A2(top_AND_M35_U1_t_reg[7]), .ZN(
        top_AND_M35_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M35_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M35_U1_OperationInst_q[5]), .A2(
        top_AND_M35_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_294) );
  OR2_X1 top_AND_M35_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M35_U1_OperationInst_q[4]), .A2(
        top_AND_M35_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M35_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M35_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M35_U1_OperationInst_q[7]), .A2(
        top_AND_M35_U1_OperationInst_q[6]), .ZN(
        top_AND_M35_U1_OperationInst_orInst2_n5) );
  OR2_X1 top_XOR_M36_U1_xorInst_U5 ( .A1(top_XOR_M36_U1_xorInst_n12), .A2(
        top_XOR_M36_U1_xorInst_n11), .ZN(top_M36) );
  INV_X1 top_XOR_M36_U1_xorInst_U4 ( .A(top_XOR_M36_U1_xorInst_n10), .ZN(
        top_XOR_M36_U1_xorInst_n11) );
  OR2_X1 top_XOR_M36_U1_xorInst_U3 ( .A1(top_XOR_M36_U1_xorInst_n9), .A2(
        top_M24), .ZN(top_XOR_M36_U1_xorInst_n10) );
  AND2_X1 top_XOR_M36_U1_xorInst_U2 ( .A1(top_M24), .A2(
        top_XOR_M36_U1_xorInst_n9), .ZN(top_XOR_M36_U1_xorInst_n12) );
  INV_X1 top_XOR_M36_U1_xorInst_U1 ( .A(Fresh[9]), .ZN(
        top_XOR_M36_U1_xorInst_n9) );
  AND2_X1 top_XOR_M36_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_271), .A2(
        top_new_AGEMA_signal_278), .ZN(top_XOR_M36_U1_w[0]) );
  AND2_X1 top_XOR_M36_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_272), .A2(
        top_new_AGEMA_signal_277), .ZN(top_XOR_M36_U1_w[1]) );
  AND2_X1 top_XOR_M36_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_272), .A2(
        top_new_AGEMA_signal_278), .ZN(top_XOR_M36_U1_w[2]) );
  AND2_X1 top_XOR_M36_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_271), .A2(
        top_new_AGEMA_signal_277), .ZN(top_XOR_M36_U1_w[3]) );
  OR2_X1 top_XOR_M36_U1_orInst1_U1 ( .A1(top_XOR_M36_U1_w[0]), .A2(
        top_XOR_M36_U1_w[1]), .ZN(top_new_AGEMA_signal_295) );
  OR2_X1 top_XOR_M36_U1_orInst2_U1 ( .A1(top_XOR_M36_U1_w[2]), .A2(
        top_XOR_M36_U1_w[3]), .ZN(top_new_AGEMA_signal_296) );
  OR2_X1 top_XOR_M37_U1_xorInst_U5 ( .A1(top_XOR_M37_U1_xorInst_n12), .A2(
        top_XOR_M37_U1_xorInst_n11), .ZN(top_M37) );
  INV_X1 top_XOR_M37_U1_xorInst_U4 ( .A(top_XOR_M37_U1_xorInst_n10), .ZN(
        top_XOR_M37_U1_xorInst_n11) );
  OR2_X1 top_XOR_M37_U1_xorInst_U3 ( .A1(top_XOR_M37_U1_xorInst_n9), .A2(
        top_M21), .ZN(top_XOR_M37_U1_xorInst_n10) );
  AND2_X1 top_XOR_M37_U1_xorInst_U2 ( .A1(top_M21), .A2(
        top_XOR_M37_U1_xorInst_n9), .ZN(top_XOR_M37_U1_xorInst_n12) );
  INV_X1 top_XOR_M37_U1_xorInst_U1 ( .A(Fresh[10]), .ZN(
        top_XOR_M37_U1_xorInst_n9) );
  AND2_X1 top_XOR_M37_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_287), .A2(
        top_new_AGEMA_signal_266), .ZN(top_XOR_M37_U1_w[0]) );
  AND2_X1 top_XOR_M37_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_288), .A2(
        top_new_AGEMA_signal_265), .ZN(top_XOR_M37_U1_w[1]) );
  AND2_X1 top_XOR_M37_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_288), .A2(
        top_new_AGEMA_signal_266), .ZN(top_XOR_M37_U1_w[2]) );
  AND2_X1 top_XOR_M37_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_287), .A2(
        top_new_AGEMA_signal_265), .ZN(top_XOR_M37_U1_w[3]) );
  OR2_X1 top_XOR_M37_U1_orInst1_U1 ( .A1(top_XOR_M37_U1_w[0]), .A2(
        top_XOR_M37_U1_w[1]), .ZN(top_new_AGEMA_signal_297) );
  OR2_X1 top_XOR_M37_U1_orInst2_U1 ( .A1(top_XOR_M37_U1_w[2]), .A2(
        top_XOR_M37_U1_w[3]), .ZN(top_new_AGEMA_signal_298) );
  OR2_X1 top_XOR_M38_U1_xorInst_U5 ( .A1(top_XOR_M38_U1_xorInst_n12), .A2(
        top_XOR_M38_U1_xorInst_n11), .ZN(top_M38) );
  INV_X1 top_XOR_M38_U1_xorInst_U4 ( .A(top_XOR_M38_U1_xorInst_n10), .ZN(
        top_XOR_M38_U1_xorInst_n11) );
  OR2_X1 top_XOR_M38_U1_xorInst_U3 ( .A1(top_XOR_M38_U1_xorInst_n9), .A2(
        Fresh[13]), .ZN(top_XOR_M38_U1_xorInst_n10) );
  AND2_X1 top_XOR_M38_U1_xorInst_U2 ( .A1(Fresh[13]), .A2(
        top_XOR_M38_U1_xorInst_n9), .ZN(top_XOR_M38_U1_xorInst_n12) );
  INV_X1 top_XOR_M38_U1_xorInst_U1 ( .A(top_M33), .ZN(
        top_XOR_M38_U1_xorInst_n9) );
  AND2_X1 top_XOR_M38_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_285), .A2(
        top_new_AGEMA_signal_292), .ZN(top_XOR_M38_U1_w[0]) );
  AND2_X1 top_XOR_M38_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_286), .A2(
        top_new_AGEMA_signal_291), .ZN(top_XOR_M38_U1_w[1]) );
  AND2_X1 top_XOR_M38_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_286), .A2(
        top_new_AGEMA_signal_292), .ZN(top_XOR_M38_U1_w[2]) );
  AND2_X1 top_XOR_M38_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_285), .A2(
        top_new_AGEMA_signal_291), .ZN(top_XOR_M38_U1_w[3]) );
  OR2_X1 top_XOR_M38_U1_orInst1_U1 ( .A1(top_XOR_M38_U1_w[0]), .A2(
        top_XOR_M38_U1_w[1]), .ZN(top_new_AGEMA_signal_299) );
  OR2_X1 top_XOR_M38_U1_orInst2_U1 ( .A1(top_XOR_M38_U1_w[2]), .A2(
        top_XOR_M38_U1_w[3]), .ZN(top_new_AGEMA_signal_300) );
  OR2_X1 top_XOR_M39_U1_xorInst_U5 ( .A1(top_XOR_M39_U1_xorInst_n12), .A2(
        top_XOR_M39_U1_xorInst_n11), .ZN(top_M39) );
  INV_X1 top_XOR_M39_U1_xorInst_U4 ( .A(top_XOR_M39_U1_xorInst_n10), .ZN(
        top_XOR_M39_U1_xorInst_n11) );
  OR2_X1 top_XOR_M39_U1_xorInst_U3 ( .A1(top_XOR_M39_U1_xorInst_n9), .A2(
        top_M23), .ZN(top_XOR_M39_U1_xorInst_n10) );
  AND2_X1 top_XOR_M39_U1_xorInst_U2 ( .A1(top_M23), .A2(
        top_XOR_M39_U1_xorInst_n9), .ZN(top_XOR_M39_U1_xorInst_n12) );
  INV_X1 top_XOR_M39_U1_xorInst_U1 ( .A(Fresh[11]), .ZN(
        top_XOR_M39_U1_xorInst_n9) );
  AND2_X1 top_XOR_M39_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_289), .A2(
        top_new_AGEMA_signal_270), .ZN(top_XOR_M39_U1_w[0]) );
  AND2_X1 top_XOR_M39_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_290), .A2(
        top_new_AGEMA_signal_269), .ZN(top_XOR_M39_U1_w[1]) );
  AND2_X1 top_XOR_M39_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_290), .A2(
        top_new_AGEMA_signal_270), .ZN(top_XOR_M39_U1_w[2]) );
  AND2_X1 top_XOR_M39_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_289), .A2(
        top_new_AGEMA_signal_269), .ZN(top_XOR_M39_U1_w[3]) );
  OR2_X1 top_XOR_M39_U1_orInst1_U1 ( .A1(top_XOR_M39_U1_w[0]), .A2(
        top_XOR_M39_U1_w[1]), .ZN(top_new_AGEMA_signal_301) );
  OR2_X1 top_XOR_M39_U1_orInst2_U1 ( .A1(top_XOR_M39_U1_w[2]), .A2(
        top_XOR_M39_U1_w[3]), .ZN(top_new_AGEMA_signal_302) );
  OR2_X1 top_XOR_M40_U1_xorInst_U5 ( .A1(top_XOR_M40_U1_xorInst_n12), .A2(
        top_XOR_M40_U1_xorInst_n11), .ZN(top_M40) );
  INV_X1 top_XOR_M40_U1_xorInst_U4 ( .A(top_XOR_M40_U1_xorInst_n10), .ZN(
        top_XOR_M40_U1_xorInst_n11) );
  OR2_X1 top_XOR_M40_U1_xorInst_U3 ( .A1(top_XOR_M40_U1_xorInst_n9), .A2(
        Fresh[15]), .ZN(top_XOR_M40_U1_xorInst_n10) );
  AND2_X1 top_XOR_M40_U1_xorInst_U2 ( .A1(Fresh[15]), .A2(
        top_XOR_M40_U1_xorInst_n9), .ZN(top_XOR_M40_U1_xorInst_n12) );
  INV_X1 top_XOR_M40_U1_xorInst_U1 ( .A(top_M36), .ZN(
        top_XOR_M40_U1_xorInst_n9) );
  AND2_X1 top_XOR_M40_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_295), .A2(
        top_new_AGEMA_signal_294), .ZN(top_XOR_M40_U1_w[0]) );
  AND2_X1 top_XOR_M40_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_296), .A2(
        top_new_AGEMA_signal_293), .ZN(top_XOR_M40_U1_w[1]) );
  AND2_X1 top_XOR_M40_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_296), .A2(
        top_new_AGEMA_signal_294), .ZN(top_XOR_M40_U1_w[2]) );
  AND2_X1 top_XOR_M40_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_295), .A2(
        top_new_AGEMA_signal_293), .ZN(top_XOR_M40_U1_w[3]) );
  OR2_X1 top_XOR_M40_U1_orInst1_U1 ( .A1(top_XOR_M40_U1_w[0]), .A2(
        top_XOR_M40_U1_w[1]), .ZN(top_new_AGEMA_signal_303) );
  OR2_X1 top_XOR_M40_U1_orInst2_U1 ( .A1(top_XOR_M40_U1_w[2]), .A2(
        top_XOR_M40_U1_w[3]), .ZN(top_new_AGEMA_signal_304) );
  OR2_X1 top_XOR_M41_U1_xorInst_U5 ( .A1(top_XOR_M41_U1_xorInst_n12), .A2(
        top_XOR_M41_U1_xorInst_n11), .ZN(top_M41) );
  INV_X1 top_XOR_M41_U1_xorInst_U4 ( .A(top_XOR_M41_U1_xorInst_n10), .ZN(
        top_XOR_M41_U1_xorInst_n11) );
  OR2_X1 top_XOR_M41_U1_xorInst_U3 ( .A1(top_XOR_M41_U1_xorInst_n9), .A2(
        top_M38), .ZN(top_XOR_M41_U1_xorInst_n10) );
  AND2_X1 top_XOR_M41_U1_xorInst_U2 ( .A1(top_M38), .A2(
        top_XOR_M41_U1_xorInst_n9), .ZN(top_XOR_M41_U1_xorInst_n12) );
  INV_X1 top_XOR_M41_U1_xorInst_U1 ( .A(top_M40), .ZN(
        top_XOR_M41_U1_xorInst_n9) );
  AND2_X1 top_XOR_M41_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_303), .A2(
        top_new_AGEMA_signal_300), .ZN(top_XOR_M41_U1_w[0]) );
  AND2_X1 top_XOR_M41_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_304), .A2(
        top_new_AGEMA_signal_299), .ZN(top_XOR_M41_U1_w[1]) );
  AND2_X1 top_XOR_M41_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_304), .A2(
        top_new_AGEMA_signal_300), .ZN(top_XOR_M41_U1_w[2]) );
  AND2_X1 top_XOR_M41_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_303), .A2(
        top_new_AGEMA_signal_299), .ZN(top_XOR_M41_U1_w[3]) );
  OR2_X1 top_XOR_M41_U1_orInst1_U1 ( .A1(top_XOR_M41_U1_w[0]), .A2(
        top_XOR_M41_U1_w[1]), .ZN(top_new_AGEMA_signal_305) );
  OR2_X1 top_XOR_M41_U1_orInst2_U1 ( .A1(top_XOR_M41_U1_w[2]), .A2(
        top_XOR_M41_U1_w[3]), .ZN(top_new_AGEMA_signal_306) );
  OR2_X1 top_XOR_M42_U1_xorInst_U5 ( .A1(top_XOR_M42_U1_xorInst_n12), .A2(
        top_XOR_M42_U1_xorInst_n11), .ZN(top_M42) );
  INV_X1 top_XOR_M42_U1_xorInst_U4 ( .A(top_XOR_M42_U1_xorInst_n10), .ZN(
        top_XOR_M42_U1_xorInst_n11) );
  OR2_X1 top_XOR_M42_U1_xorInst_U3 ( .A1(top_XOR_M42_U1_xorInst_n9), .A2(
        top_M37), .ZN(top_XOR_M42_U1_xorInst_n10) );
  AND2_X1 top_XOR_M42_U1_xorInst_U2 ( .A1(top_M37), .A2(
        top_XOR_M42_U1_xorInst_n9), .ZN(top_XOR_M42_U1_xorInst_n12) );
  INV_X1 top_XOR_M42_U1_xorInst_U1 ( .A(top_M39), .ZN(
        top_XOR_M42_U1_xorInst_n9) );
  AND2_X1 top_XOR_M42_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_301), .A2(
        top_new_AGEMA_signal_298), .ZN(top_XOR_M42_U1_w[0]) );
  AND2_X1 top_XOR_M42_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_302), .A2(
        top_new_AGEMA_signal_297), .ZN(top_XOR_M42_U1_w[1]) );
  AND2_X1 top_XOR_M42_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_302), .A2(
        top_new_AGEMA_signal_298), .ZN(top_XOR_M42_U1_w[2]) );
  AND2_X1 top_XOR_M42_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_301), .A2(
        top_new_AGEMA_signal_297), .ZN(top_XOR_M42_U1_w[3]) );
  OR2_X1 top_XOR_M42_U1_orInst1_U1 ( .A1(top_XOR_M42_U1_w[0]), .A2(
        top_XOR_M42_U1_w[1]), .ZN(top_new_AGEMA_signal_307) );
  OR2_X1 top_XOR_M42_U1_orInst2_U1 ( .A1(top_XOR_M42_U1_w[2]), .A2(
        top_XOR_M42_U1_w[3]), .ZN(top_new_AGEMA_signal_308) );
  OR2_X1 top_XOR_M43_U1_xorInst_U5 ( .A1(top_XOR_M43_U1_xorInst_n12), .A2(
        top_XOR_M43_U1_xorInst_n11), .ZN(top_M43) );
  INV_X1 top_XOR_M43_U1_xorInst_U4 ( .A(top_XOR_M43_U1_xorInst_n10), .ZN(
        top_XOR_M43_U1_xorInst_n11) );
  OR2_X1 top_XOR_M43_U1_xorInst_U3 ( .A1(top_XOR_M43_U1_xorInst_n9), .A2(
        top_M37), .ZN(top_XOR_M43_U1_xorInst_n10) );
  AND2_X1 top_XOR_M43_U1_xorInst_U2 ( .A1(top_M37), .A2(
        top_XOR_M43_U1_xorInst_n9), .ZN(top_XOR_M43_U1_xorInst_n12) );
  INV_X1 top_XOR_M43_U1_xorInst_U1 ( .A(top_M38), .ZN(
        top_XOR_M43_U1_xorInst_n9) );
  AND2_X1 top_XOR_M43_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_299), .A2(
        top_new_AGEMA_signal_298), .ZN(top_XOR_M43_U1_w[0]) );
  AND2_X1 top_XOR_M43_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_300), .A2(
        top_new_AGEMA_signal_297), .ZN(top_XOR_M43_U1_w[1]) );
  AND2_X1 top_XOR_M43_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_300), .A2(
        top_new_AGEMA_signal_298), .ZN(top_XOR_M43_U1_w[2]) );
  AND2_X1 top_XOR_M43_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_299), .A2(
        top_new_AGEMA_signal_297), .ZN(top_XOR_M43_U1_w[3]) );
  OR2_X1 top_XOR_M43_U1_orInst1_U1 ( .A1(top_XOR_M43_U1_w[0]), .A2(
        top_XOR_M43_U1_w[1]), .ZN(top_new_AGEMA_signal_309) );
  OR2_X1 top_XOR_M43_U1_orInst2_U1 ( .A1(top_XOR_M43_U1_w[2]), .A2(
        top_XOR_M43_U1_w[3]), .ZN(top_new_AGEMA_signal_310) );
  OR2_X1 top_XOR_M44_U1_xorInst_U5 ( .A1(top_XOR_M44_U1_xorInst_n12), .A2(
        top_XOR_M44_U1_xorInst_n11), .ZN(top_M44) );
  INV_X1 top_XOR_M44_U1_xorInst_U4 ( .A(top_XOR_M44_U1_xorInst_n10), .ZN(
        top_XOR_M44_U1_xorInst_n11) );
  OR2_X1 top_XOR_M44_U1_xorInst_U3 ( .A1(top_XOR_M44_U1_xorInst_n9), .A2(
        top_M39), .ZN(top_XOR_M44_U1_xorInst_n10) );
  AND2_X1 top_XOR_M44_U1_xorInst_U2 ( .A1(top_M39), .A2(
        top_XOR_M44_U1_xorInst_n9), .ZN(top_XOR_M44_U1_xorInst_n12) );
  INV_X1 top_XOR_M44_U1_xorInst_U1 ( .A(top_M40), .ZN(
        top_XOR_M44_U1_xorInst_n9) );
  AND2_X1 top_XOR_M44_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_303), .A2(
        top_new_AGEMA_signal_302), .ZN(top_XOR_M44_U1_w[0]) );
  AND2_X1 top_XOR_M44_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_304), .A2(
        top_new_AGEMA_signal_301), .ZN(top_XOR_M44_U1_w[1]) );
  AND2_X1 top_XOR_M44_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_304), .A2(
        top_new_AGEMA_signal_302), .ZN(top_XOR_M44_U1_w[2]) );
  AND2_X1 top_XOR_M44_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_303), .A2(
        top_new_AGEMA_signal_301), .ZN(top_XOR_M44_U1_w[3]) );
  OR2_X1 top_XOR_M44_U1_orInst1_U1 ( .A1(top_XOR_M44_U1_w[0]), .A2(
        top_XOR_M44_U1_w[1]), .ZN(top_new_AGEMA_signal_311) );
  OR2_X1 top_XOR_M44_U1_orInst2_U1 ( .A1(top_XOR_M44_U1_w[2]), .A2(
        top_XOR_M44_U1_w[3]), .ZN(top_new_AGEMA_signal_312) );
  OR2_X1 top_XOR_M45_U1_xorInst_U5 ( .A1(top_XOR_M45_U1_xorInst_n12), .A2(
        top_XOR_M45_U1_xorInst_n11), .ZN(top_M45) );
  INV_X1 top_XOR_M45_U1_xorInst_U4 ( .A(top_XOR_M45_U1_xorInst_n10), .ZN(
        top_XOR_M45_U1_xorInst_n11) );
  OR2_X1 top_XOR_M45_U1_xorInst_U3 ( .A1(top_XOR_M45_U1_xorInst_n9), .A2(
        top_M42), .ZN(top_XOR_M45_U1_xorInst_n10) );
  AND2_X1 top_XOR_M45_U1_xorInst_U2 ( .A1(top_M42), .A2(
        top_XOR_M45_U1_xorInst_n9), .ZN(top_XOR_M45_U1_xorInst_n12) );
  INV_X1 top_XOR_M45_U1_xorInst_U1 ( .A(top_M41), .ZN(
        top_XOR_M45_U1_xorInst_n9) );
  AND2_X1 top_XOR_M45_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_305), .A2(
        top_new_AGEMA_signal_308), .ZN(top_XOR_M45_U1_w[0]) );
  AND2_X1 top_XOR_M45_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_306), .A2(
        top_new_AGEMA_signal_307), .ZN(top_XOR_M45_U1_w[1]) );
  AND2_X1 top_XOR_M45_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_306), .A2(
        top_new_AGEMA_signal_308), .ZN(top_XOR_M45_U1_w[2]) );
  AND2_X1 top_XOR_M45_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_305), .A2(
        top_new_AGEMA_signal_307), .ZN(top_XOR_M45_U1_w[3]) );
  OR2_X1 top_XOR_M45_U1_orInst1_U1 ( .A1(top_XOR_M45_U1_w[0]), .A2(
        top_XOR_M45_U1_w[1]), .ZN(top_new_AGEMA_signal_329) );
  OR2_X1 top_XOR_M45_U1_orInst2_U1 ( .A1(top_XOR_M45_U1_w[2]), .A2(
        top_XOR_M45_U1_w[3]), .ZN(top_new_AGEMA_signal_330) );
  INV_X1 top_AND_M46_U1_nonlinearInst_U26 ( .A(top_AND_M46_U1_t[3]), .ZN(
        top_AND_M46_U1_t[7]) );
  OR2_X1 top_AND_M46_U1_nonlinearInst_U25 ( .A1(
        top_AND_M46_U1_nonlinearInst_n64), .A2(
        top_AND_M46_U1_nonlinearInst_n63), .ZN(top_AND_M46_U1_t[3]) );
  INV_X1 top_AND_M46_U1_nonlinearInst_U24 ( .A(
        top_AND_M46_U1_nonlinearInst_n62), .ZN(
        top_AND_M46_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M46_U1_nonlinearInst_U23 ( .A1(
        top_AND_M46_U1_nonlinearInst_n61), .A2(Fresh[16]), .ZN(
        top_AND_M46_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M46_U1_nonlinearInst_U22 ( .A1(Fresh[16]), .A2(
        top_AND_M46_U1_nonlinearInst_n61), .ZN(
        top_AND_M46_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M46_U1_nonlinearInst_U21 ( .A1(top_M44), .A2(top_T6), .ZN(
        top_AND_M46_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M46_U1_nonlinearInst_U20 ( .A(top_AND_M46_U1_t[2]), .ZN(
        top_AND_M46_U1_t[6]) );
  OR2_X1 top_AND_M46_U1_nonlinearInst_U19 ( .A1(
        top_AND_M46_U1_nonlinearInst_n60), .A2(
        top_AND_M46_U1_nonlinearInst_n59), .ZN(top_AND_M46_U1_t[2]) );
  INV_X1 top_AND_M46_U1_nonlinearInst_U18 ( .A(
        top_AND_M46_U1_nonlinearInst_n58), .ZN(
        top_AND_M46_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M46_U1_nonlinearInst_U17 ( .A1(
        top_AND_M46_U1_nonlinearInst_n57), .A2(Fresh[16]), .ZN(
        top_AND_M46_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M46_U1_nonlinearInst_U16 ( .A1(Fresh[16]), .A2(
        top_AND_M46_U1_nonlinearInst_n57), .ZN(
        top_AND_M46_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M46_U1_nonlinearInst_U15 ( .A1(
        top_AND_M46_U1_nonlinearInst_n56), .A2(top_M44), .ZN(
        top_AND_M46_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M46_U1_nonlinearInst_U14 ( .A(top_AND_M46_U1_t[1]), .ZN(
        top_AND_M46_U1_t[5]) );
  OR2_X1 top_AND_M46_U1_nonlinearInst_U13 ( .A1(
        top_AND_M46_U1_nonlinearInst_n55), .A2(
        top_AND_M46_U1_nonlinearInst_n54), .ZN(top_AND_M46_U1_t[1]) );
  AND2_X1 top_AND_M46_U1_nonlinearInst_U12 ( .A1(
        top_AND_M46_U1_nonlinearInst_n53), .A2(
        top_AND_M46_U1_nonlinearInst_n52), .ZN(
        top_AND_M46_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M46_U1_nonlinearInst_U11 ( .A(
        top_AND_M46_U1_nonlinearInst_n51), .ZN(
        top_AND_M46_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M46_U1_nonlinearInst_U10 ( .A1(
        top_AND_M46_U1_nonlinearInst_n52), .A2(
        top_AND_M46_U1_nonlinearInst_n53), .ZN(
        top_AND_M46_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M46_U1_nonlinearInst_U9 ( .A1(top_M44), .A2(
        top_AND_M46_U1_nonlinearInst_n56), .ZN(
        top_AND_M46_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M46_U1_nonlinearInst_U8 ( .A(top_T6), .ZN(
        top_AND_M46_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M46_U1_nonlinearInst_U7 ( .A(top_AND_M46_U1_t[0]), .ZN(
        top_AND_M46_U1_t[4]) );
  OR2_X1 top_AND_M46_U1_nonlinearInst_U6 ( .A1(
        top_AND_M46_U1_nonlinearInst_n50), .A2(
        top_AND_M46_U1_nonlinearInst_n49), .ZN(top_AND_M46_U1_t[0]) );
  AND2_X1 top_AND_M46_U1_nonlinearInst_U5 ( .A1(
        top_AND_M46_U1_nonlinearInst_n48), .A2(
        top_AND_M46_U1_nonlinearInst_n52), .ZN(
        top_AND_M46_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M46_U1_nonlinearInst_U4 ( .A(top_AND_M46_U1_nonlinearInst_n47), .ZN(top_AND_M46_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M46_U1_nonlinearInst_U3 ( .A1(
        top_AND_M46_U1_nonlinearInst_n52), .A2(
        top_AND_M46_U1_nonlinearInst_n48), .ZN(
        top_AND_M46_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M46_U1_nonlinearInst_U2 ( .A1(top_M44), .A2(top_T6), .ZN(
        top_AND_M46_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M46_U1_nonlinearInst_U1 ( .A(Fresh[16]), .ZN(
        top_AND_M46_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M46_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M46_U1_t[0]), .A2(
        top_AND_M46_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M46_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M46_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M46_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M46_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M46_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M46_U1_t_reg[0]) );
  AND2_X1 top_AND_M46_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M46_U1_t[1]), .A2(
        top_AND_M46_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M46_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M46_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M46_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M46_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M46_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M46_U1_t_reg[1]) );
  AND2_X1 top_AND_M46_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M46_U1_t[2]), .A2(
        top_AND_M46_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M46_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M46_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M46_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M46_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M46_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M46_U1_t_reg[2]) );
  AND2_X1 top_AND_M46_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M46_U1_t[3]), .A2(
        top_AND_M46_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M46_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M46_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M46_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M46_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M46_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M46_U1_t_reg[3]) );
  AND2_X1 top_AND_M46_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M46_U1_t[4]), .A2(
        top_AND_M46_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M46_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M46_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M46_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M46_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M46_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M46_U1_t_reg[4]) );
  AND2_X1 top_AND_M46_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M46_U1_t[5]), .A2(
        top_AND_M46_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M46_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M46_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M46_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M46_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M46_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M46_U1_t_reg[5]) );
  AND2_X1 top_AND_M46_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M46_U1_t[6]), .A2(
        top_AND_M46_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M46_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M46_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M46_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M46_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M46_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M46_U1_t_reg[6]) );
  AND2_X1 top_AND_M46_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M46_U1_t[7]), .A2(
        top_AND_M46_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M46_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M46_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M46_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M46_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M46_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M46_U1_t_reg[7]) );
  AND2_X1 top_AND_M46_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_192), .A2(
        top_AND_M46_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M46_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M46_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_312), .A2(top_AND_M46_U1_t_reg[0]), .ZN(
        top_AND_M46_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M46_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_191), .A2(
        top_AND_M46_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M46_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M46_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_312), .A2(top_AND_M46_U1_t_reg[1]), .ZN(
        top_AND_M46_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M46_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_192), .A2(
        top_AND_M46_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M46_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M46_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_311), .A2(top_AND_M46_U1_t_reg[2]), .ZN(
        top_AND_M46_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M46_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_191), .A2(
        top_AND_M46_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M46_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M46_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_311), .A2(top_AND_M46_U1_t_reg[3]), .ZN(
        top_AND_M46_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M46_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M46_U1_OperationInst_q[1]), .A2(
        top_AND_M46_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_331) );
  OR2_X1 top_AND_M46_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M46_U1_OperationInst_q[0]), .A2(
        top_AND_M46_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M46_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M46_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M46_U1_OperationInst_q[3]), .A2(
        top_AND_M46_U1_OperationInst_q[2]), .ZN(
        top_AND_M46_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M46_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_192), .A2(
        top_AND_M46_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M46_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M46_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_312), .A2(top_AND_M46_U1_t_reg[4]), .ZN(
        top_AND_M46_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M46_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_191), .A2(
        top_AND_M46_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M46_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M46_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_312), .A2(top_AND_M46_U1_t_reg[5]), .ZN(
        top_AND_M46_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M46_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_192), .A2(
        top_AND_M46_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M46_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M46_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_311), .A2(top_AND_M46_U1_t_reg[6]), .ZN(
        top_AND_M46_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M46_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_191), .A2(
        top_AND_M46_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M46_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M46_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_311), .A2(top_AND_M46_U1_t_reg[7]), .ZN(
        top_AND_M46_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M46_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M46_U1_OperationInst_q[5]), .A2(
        top_AND_M46_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_332) );
  OR2_X1 top_AND_M46_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M46_U1_OperationInst_q[4]), .A2(
        top_AND_M46_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M46_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M46_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M46_U1_OperationInst_q[7]), .A2(
        top_AND_M46_U1_OperationInst_q[6]), .ZN(
        top_AND_M46_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M47_U1_nonlinearInst_U26 ( .A(top_AND_M47_U1_t[3]), .ZN(
        top_AND_M47_U1_t[7]) );
  OR2_X1 top_AND_M47_U1_nonlinearInst_U25 ( .A1(
        top_AND_M47_U1_nonlinearInst_n64), .A2(
        top_AND_M47_U1_nonlinearInst_n63), .ZN(top_AND_M47_U1_t[3]) );
  INV_X1 top_AND_M47_U1_nonlinearInst_U24 ( .A(
        top_AND_M47_U1_nonlinearInst_n62), .ZN(
        top_AND_M47_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M47_U1_nonlinearInst_U23 ( .A1(
        top_AND_M47_U1_nonlinearInst_n61), .A2(Fresh[17]), .ZN(
        top_AND_M47_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M47_U1_nonlinearInst_U22 ( .A1(Fresh[17]), .A2(
        top_AND_M47_U1_nonlinearInst_n61), .ZN(
        top_AND_M47_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M47_U1_nonlinearInst_U21 ( .A1(top_M40), .A2(top_T8), .ZN(
        top_AND_M47_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M47_U1_nonlinearInst_U20 ( .A(top_AND_M47_U1_t[2]), .ZN(
        top_AND_M47_U1_t[6]) );
  OR2_X1 top_AND_M47_U1_nonlinearInst_U19 ( .A1(
        top_AND_M47_U1_nonlinearInst_n60), .A2(
        top_AND_M47_U1_nonlinearInst_n59), .ZN(top_AND_M47_U1_t[2]) );
  INV_X1 top_AND_M47_U1_nonlinearInst_U18 ( .A(
        top_AND_M47_U1_nonlinearInst_n58), .ZN(
        top_AND_M47_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M47_U1_nonlinearInst_U17 ( .A1(
        top_AND_M47_U1_nonlinearInst_n57), .A2(Fresh[17]), .ZN(
        top_AND_M47_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M47_U1_nonlinearInst_U16 ( .A1(Fresh[17]), .A2(
        top_AND_M47_U1_nonlinearInst_n57), .ZN(
        top_AND_M47_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M47_U1_nonlinearInst_U15 ( .A1(
        top_AND_M47_U1_nonlinearInst_n56), .A2(top_M40), .ZN(
        top_AND_M47_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M47_U1_nonlinearInst_U14 ( .A(top_AND_M47_U1_t[1]), .ZN(
        top_AND_M47_U1_t[5]) );
  OR2_X1 top_AND_M47_U1_nonlinearInst_U13 ( .A1(
        top_AND_M47_U1_nonlinearInst_n55), .A2(
        top_AND_M47_U1_nonlinearInst_n54), .ZN(top_AND_M47_U1_t[1]) );
  AND2_X1 top_AND_M47_U1_nonlinearInst_U12 ( .A1(
        top_AND_M47_U1_nonlinearInst_n53), .A2(
        top_AND_M47_U1_nonlinearInst_n52), .ZN(
        top_AND_M47_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M47_U1_nonlinearInst_U11 ( .A(
        top_AND_M47_U1_nonlinearInst_n51), .ZN(
        top_AND_M47_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M47_U1_nonlinearInst_U10 ( .A1(
        top_AND_M47_U1_nonlinearInst_n52), .A2(
        top_AND_M47_U1_nonlinearInst_n53), .ZN(
        top_AND_M47_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M47_U1_nonlinearInst_U9 ( .A1(top_M40), .A2(
        top_AND_M47_U1_nonlinearInst_n56), .ZN(
        top_AND_M47_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M47_U1_nonlinearInst_U8 ( .A(top_T8), .ZN(
        top_AND_M47_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M47_U1_nonlinearInst_U7 ( .A(top_AND_M47_U1_t[0]), .ZN(
        top_AND_M47_U1_t[4]) );
  OR2_X1 top_AND_M47_U1_nonlinearInst_U6 ( .A1(
        top_AND_M47_U1_nonlinearInst_n50), .A2(
        top_AND_M47_U1_nonlinearInst_n49), .ZN(top_AND_M47_U1_t[0]) );
  AND2_X1 top_AND_M47_U1_nonlinearInst_U5 ( .A1(
        top_AND_M47_U1_nonlinearInst_n48), .A2(
        top_AND_M47_U1_nonlinearInst_n52), .ZN(
        top_AND_M47_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M47_U1_nonlinearInst_U4 ( .A(top_AND_M47_U1_nonlinearInst_n47), .ZN(top_AND_M47_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M47_U1_nonlinearInst_U3 ( .A1(
        top_AND_M47_U1_nonlinearInst_n52), .A2(
        top_AND_M47_U1_nonlinearInst_n48), .ZN(
        top_AND_M47_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M47_U1_nonlinearInst_U2 ( .A1(top_M40), .A2(top_T8), .ZN(
        top_AND_M47_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M47_U1_nonlinearInst_U1 ( .A(Fresh[17]), .ZN(
        top_AND_M47_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M47_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M47_U1_t[0]), .A2(
        top_AND_M47_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M47_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M47_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M47_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M47_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M47_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M47_U1_t_reg[0]) );
  AND2_X1 top_AND_M47_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M47_U1_t[1]), .A2(
        top_AND_M47_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M47_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M47_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M47_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M47_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M47_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M47_U1_t_reg[1]) );
  AND2_X1 top_AND_M47_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M47_U1_t[2]), .A2(
        top_AND_M47_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M47_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M47_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M47_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M47_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M47_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M47_U1_t_reg[2]) );
  AND2_X1 top_AND_M47_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M47_U1_t[3]), .A2(
        top_AND_M47_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M47_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M47_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M47_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M47_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M47_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M47_U1_t_reg[3]) );
  AND2_X1 top_AND_M47_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M47_U1_t[4]), .A2(
        top_AND_M47_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M47_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M47_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M47_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M47_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M47_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M47_U1_t_reg[4]) );
  AND2_X1 top_AND_M47_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M47_U1_t[5]), .A2(
        top_AND_M47_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M47_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M47_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M47_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M47_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M47_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M47_U1_t_reg[5]) );
  AND2_X1 top_AND_M47_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M47_U1_t[6]), .A2(
        top_AND_M47_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M47_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M47_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M47_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M47_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M47_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M47_U1_t_reg[6]) );
  AND2_X1 top_AND_M47_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M47_U1_t[7]), .A2(
        top_AND_M47_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M47_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M47_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M47_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M47_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M47_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M47_U1_t_reg[7]) );
  AND2_X1 top_AND_M47_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_208), .A2(
        top_AND_M47_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M47_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M47_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_304), .A2(top_AND_M47_U1_t_reg[0]), .ZN(
        top_AND_M47_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M47_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_207), .A2(
        top_AND_M47_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M47_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M47_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_304), .A2(top_AND_M47_U1_t_reg[1]), .ZN(
        top_AND_M47_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M47_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_208), .A2(
        top_AND_M47_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M47_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M47_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_303), .A2(top_AND_M47_U1_t_reg[2]), .ZN(
        top_AND_M47_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M47_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_207), .A2(
        top_AND_M47_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M47_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M47_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_303), .A2(top_AND_M47_U1_t_reg[3]), .ZN(
        top_AND_M47_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M47_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M47_U1_OperationInst_q[1]), .A2(
        top_AND_M47_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_313) );
  OR2_X1 top_AND_M47_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M47_U1_OperationInst_q[0]), .A2(
        top_AND_M47_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M47_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M47_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M47_U1_OperationInst_q[3]), .A2(
        top_AND_M47_U1_OperationInst_q[2]), .ZN(
        top_AND_M47_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M47_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_208), .A2(
        top_AND_M47_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M47_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M47_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_304), .A2(top_AND_M47_U1_t_reg[4]), .ZN(
        top_AND_M47_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M47_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_207), .A2(
        top_AND_M47_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M47_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M47_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_304), .A2(top_AND_M47_U1_t_reg[5]), .ZN(
        top_AND_M47_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M47_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_208), .A2(
        top_AND_M47_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M47_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M47_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_303), .A2(top_AND_M47_U1_t_reg[6]), .ZN(
        top_AND_M47_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M47_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_207), .A2(
        top_AND_M47_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M47_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M47_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_303), .A2(top_AND_M47_U1_t_reg[7]), .ZN(
        top_AND_M47_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M47_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M47_U1_OperationInst_q[5]), .A2(
        top_AND_M47_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_314) );
  OR2_X1 top_AND_M47_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M47_U1_OperationInst_q[4]), .A2(
        top_AND_M47_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M47_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M47_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M47_U1_OperationInst_q[7]), .A2(
        top_AND_M47_U1_OperationInst_q[6]), .ZN(
        top_AND_M47_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M48_U1_nonlinearInst_U26 ( .A(top_AND_M48_U1_t[3]), .ZN(
        top_AND_M48_U1_t[7]) );
  OR2_X1 top_AND_M48_U1_nonlinearInst_U25 ( .A1(
        top_AND_M48_U1_nonlinearInst_n64), .A2(
        top_AND_M48_U1_nonlinearInst_n63), .ZN(top_AND_M48_U1_t[3]) );
  INV_X1 top_AND_M48_U1_nonlinearInst_U24 ( .A(
        top_AND_M48_U1_nonlinearInst_n62), .ZN(
        top_AND_M48_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M48_U1_nonlinearInst_U23 ( .A1(
        top_AND_M48_U1_nonlinearInst_n61), .A2(Fresh[18]), .ZN(
        top_AND_M48_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M48_U1_nonlinearInst_U22 ( .A1(Fresh[18]), .A2(
        top_AND_M48_U1_nonlinearInst_n61), .ZN(
        top_AND_M48_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M48_U1_nonlinearInst_U21 ( .A1(top_M39), .A2(X_s0[0]), .ZN(
        top_AND_M48_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M48_U1_nonlinearInst_U20 ( .A(top_AND_M48_U1_t[2]), .ZN(
        top_AND_M48_U1_t[6]) );
  OR2_X1 top_AND_M48_U1_nonlinearInst_U19 ( .A1(
        top_AND_M48_U1_nonlinearInst_n60), .A2(
        top_AND_M48_U1_nonlinearInst_n59), .ZN(top_AND_M48_U1_t[2]) );
  INV_X1 top_AND_M48_U1_nonlinearInst_U18 ( .A(
        top_AND_M48_U1_nonlinearInst_n58), .ZN(
        top_AND_M48_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M48_U1_nonlinearInst_U17 ( .A1(
        top_AND_M48_U1_nonlinearInst_n57), .A2(Fresh[18]), .ZN(
        top_AND_M48_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M48_U1_nonlinearInst_U16 ( .A1(Fresh[18]), .A2(
        top_AND_M48_U1_nonlinearInst_n57), .ZN(
        top_AND_M48_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M48_U1_nonlinearInst_U15 ( .A1(
        top_AND_M48_U1_nonlinearInst_n56), .A2(top_M39), .ZN(
        top_AND_M48_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M48_U1_nonlinearInst_U14 ( .A(top_AND_M48_U1_t[1]), .ZN(
        top_AND_M48_U1_t[5]) );
  OR2_X1 top_AND_M48_U1_nonlinearInst_U13 ( .A1(
        top_AND_M48_U1_nonlinearInst_n55), .A2(
        top_AND_M48_U1_nonlinearInst_n54), .ZN(top_AND_M48_U1_t[1]) );
  AND2_X1 top_AND_M48_U1_nonlinearInst_U12 ( .A1(
        top_AND_M48_U1_nonlinearInst_n53), .A2(
        top_AND_M48_U1_nonlinearInst_n52), .ZN(
        top_AND_M48_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M48_U1_nonlinearInst_U11 ( .A(
        top_AND_M48_U1_nonlinearInst_n51), .ZN(
        top_AND_M48_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M48_U1_nonlinearInst_U10 ( .A1(
        top_AND_M48_U1_nonlinearInst_n52), .A2(
        top_AND_M48_U1_nonlinearInst_n53), .ZN(
        top_AND_M48_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M48_U1_nonlinearInst_U9 ( .A1(top_M39), .A2(
        top_AND_M48_U1_nonlinearInst_n56), .ZN(
        top_AND_M48_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M48_U1_nonlinearInst_U8 ( .A(X_s0[0]), .ZN(
        top_AND_M48_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M48_U1_nonlinearInst_U7 ( .A(top_AND_M48_U1_t[0]), .ZN(
        top_AND_M48_U1_t[4]) );
  OR2_X1 top_AND_M48_U1_nonlinearInst_U6 ( .A1(
        top_AND_M48_U1_nonlinearInst_n50), .A2(
        top_AND_M48_U1_nonlinearInst_n49), .ZN(top_AND_M48_U1_t[0]) );
  AND2_X1 top_AND_M48_U1_nonlinearInst_U5 ( .A1(
        top_AND_M48_U1_nonlinearInst_n48), .A2(
        top_AND_M48_U1_nonlinearInst_n52), .ZN(
        top_AND_M48_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M48_U1_nonlinearInst_U4 ( .A(top_AND_M48_U1_nonlinearInst_n47), .ZN(top_AND_M48_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M48_U1_nonlinearInst_U3 ( .A1(
        top_AND_M48_U1_nonlinearInst_n52), .A2(
        top_AND_M48_U1_nonlinearInst_n48), .ZN(
        top_AND_M48_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M48_U1_nonlinearInst_U2 ( .A1(top_M39), .A2(X_s0[0]), .ZN(
        top_AND_M48_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M48_U1_nonlinearInst_U1 ( .A(Fresh[18]), .ZN(
        top_AND_M48_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M48_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M48_U1_t[0]), .A2(
        top_AND_M48_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M48_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M48_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M48_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M48_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M48_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M48_U1_t_reg[0]) );
  AND2_X1 top_AND_M48_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M48_U1_t[1]), .A2(
        top_AND_M48_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M48_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M48_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M48_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M48_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M48_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M48_U1_t_reg[1]) );
  AND2_X1 top_AND_M48_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M48_U1_t[2]), .A2(
        top_AND_M48_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M48_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M48_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M48_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M48_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M48_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M48_U1_t_reg[2]) );
  AND2_X1 top_AND_M48_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M48_U1_t[3]), .A2(
        top_AND_M48_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M48_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M48_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M48_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M48_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M48_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M48_U1_t_reg[3]) );
  AND2_X1 top_AND_M48_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M48_U1_t[4]), .A2(
        top_AND_M48_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M48_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M48_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M48_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M48_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M48_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M48_U1_t_reg[4]) );
  AND2_X1 top_AND_M48_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M48_U1_t[5]), .A2(
        top_AND_M48_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M48_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M48_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M48_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M48_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M48_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M48_U1_t_reg[5]) );
  AND2_X1 top_AND_M48_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M48_U1_t[6]), .A2(
        top_AND_M48_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M48_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M48_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M48_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M48_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M48_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M48_U1_t_reg[6]) );
  AND2_X1 top_AND_M48_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M48_U1_t[7]), .A2(
        top_AND_M48_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M48_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M48_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M48_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M48_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M48_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M48_U1_t_reg[7]) );
  AND2_X1 top_AND_M48_U1_OperationInst_andInst0_U2 ( .A1(X_s1_bar[0]), .A2(
        top_AND_M48_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M48_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M48_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_302), .A2(top_AND_M48_U1_t_reg[0]), .ZN(
        top_AND_M48_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M48_U1_OperationInst_andInst1_U2 ( .A1(X_s1[0]), .A2(
        top_AND_M48_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M48_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M48_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_302), .A2(top_AND_M48_U1_t_reg[1]), .ZN(
        top_AND_M48_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M48_U1_OperationInst_andInst2_U2 ( .A1(X_s1_bar[0]), .A2(
        top_AND_M48_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M48_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M48_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_301), .A2(top_AND_M48_U1_t_reg[2]), .ZN(
        top_AND_M48_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M48_U1_OperationInst_andInst3_U2 ( .A1(X_s1[0]), .A2(
        top_AND_M48_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M48_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M48_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_301), .A2(top_AND_M48_U1_t_reg[3]), .ZN(
        top_AND_M48_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M48_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M48_U1_OperationInst_q[1]), .A2(
        top_AND_M48_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_315) );
  OR2_X1 top_AND_M48_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M48_U1_OperationInst_q[0]), .A2(
        top_AND_M48_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M48_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M48_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M48_U1_OperationInst_q[3]), .A2(
        top_AND_M48_U1_OperationInst_q[2]), .ZN(
        top_AND_M48_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M48_U1_OperationInst_andInst4_U2 ( .A1(X_s1_bar[0]), .A2(
        top_AND_M48_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M48_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M48_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_302), .A2(top_AND_M48_U1_t_reg[4]), .ZN(
        top_AND_M48_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M48_U1_OperationInst_andInst5_U2 ( .A1(X_s1[0]), .A2(
        top_AND_M48_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M48_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M48_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_302), .A2(top_AND_M48_U1_t_reg[5]), .ZN(
        top_AND_M48_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M48_U1_OperationInst_andInst6_U2 ( .A1(X_s1_bar[0]), .A2(
        top_AND_M48_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M48_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M48_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_301), .A2(top_AND_M48_U1_t_reg[6]), .ZN(
        top_AND_M48_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M48_U1_OperationInst_andInst7_U2 ( .A1(X_s1[0]), .A2(
        top_AND_M48_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M48_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M48_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_301), .A2(top_AND_M48_U1_t_reg[7]), .ZN(
        top_AND_M48_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M48_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M48_U1_OperationInst_q[5]), .A2(
        top_AND_M48_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_316) );
  OR2_X1 top_AND_M48_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M48_U1_OperationInst_q[4]), .A2(
        top_AND_M48_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M48_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M48_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M48_U1_OperationInst_q[7]), .A2(
        top_AND_M48_U1_OperationInst_q[6]), .ZN(
        top_AND_M48_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M49_U1_nonlinearInst_U26 ( .A(top_AND_M49_U1_t[3]), .ZN(
        top_AND_M49_U1_t[7]) );
  OR2_X1 top_AND_M49_U1_nonlinearInst_U25 ( .A1(
        top_AND_M49_U1_nonlinearInst_n64), .A2(
        top_AND_M49_U1_nonlinearInst_n63), .ZN(top_AND_M49_U1_t[3]) );
  INV_X1 top_AND_M49_U1_nonlinearInst_U24 ( .A(
        top_AND_M49_U1_nonlinearInst_n62), .ZN(
        top_AND_M49_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M49_U1_nonlinearInst_U23 ( .A1(
        top_AND_M49_U1_nonlinearInst_n61), .A2(Fresh[19]), .ZN(
        top_AND_M49_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M49_U1_nonlinearInst_U22 ( .A1(Fresh[19]), .A2(
        top_AND_M49_U1_nonlinearInst_n61), .ZN(
        top_AND_M49_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M49_U1_nonlinearInst_U21 ( .A1(top_M43), .A2(top_T16), .ZN(
        top_AND_M49_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M49_U1_nonlinearInst_U20 ( .A(top_AND_M49_U1_t[2]), .ZN(
        top_AND_M49_U1_t[6]) );
  OR2_X1 top_AND_M49_U1_nonlinearInst_U19 ( .A1(
        top_AND_M49_U1_nonlinearInst_n60), .A2(
        top_AND_M49_U1_nonlinearInst_n59), .ZN(top_AND_M49_U1_t[2]) );
  INV_X1 top_AND_M49_U1_nonlinearInst_U18 ( .A(
        top_AND_M49_U1_nonlinearInst_n58), .ZN(
        top_AND_M49_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M49_U1_nonlinearInst_U17 ( .A1(
        top_AND_M49_U1_nonlinearInst_n57), .A2(Fresh[19]), .ZN(
        top_AND_M49_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M49_U1_nonlinearInst_U16 ( .A1(Fresh[19]), .A2(
        top_AND_M49_U1_nonlinearInst_n57), .ZN(
        top_AND_M49_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M49_U1_nonlinearInst_U15 ( .A1(
        top_AND_M49_U1_nonlinearInst_n56), .A2(top_M43), .ZN(
        top_AND_M49_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M49_U1_nonlinearInst_U14 ( .A(top_AND_M49_U1_t[1]), .ZN(
        top_AND_M49_U1_t[5]) );
  OR2_X1 top_AND_M49_U1_nonlinearInst_U13 ( .A1(
        top_AND_M49_U1_nonlinearInst_n55), .A2(
        top_AND_M49_U1_nonlinearInst_n54), .ZN(top_AND_M49_U1_t[1]) );
  AND2_X1 top_AND_M49_U1_nonlinearInst_U12 ( .A1(
        top_AND_M49_U1_nonlinearInst_n53), .A2(
        top_AND_M49_U1_nonlinearInst_n52), .ZN(
        top_AND_M49_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M49_U1_nonlinearInst_U11 ( .A(
        top_AND_M49_U1_nonlinearInst_n51), .ZN(
        top_AND_M49_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M49_U1_nonlinearInst_U10 ( .A1(
        top_AND_M49_U1_nonlinearInst_n52), .A2(
        top_AND_M49_U1_nonlinearInst_n53), .ZN(
        top_AND_M49_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M49_U1_nonlinearInst_U9 ( .A1(top_M43), .A2(
        top_AND_M49_U1_nonlinearInst_n56), .ZN(
        top_AND_M49_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M49_U1_nonlinearInst_U8 ( .A(top_T16), .ZN(
        top_AND_M49_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M49_U1_nonlinearInst_U7 ( .A(top_AND_M49_U1_t[0]), .ZN(
        top_AND_M49_U1_t[4]) );
  OR2_X1 top_AND_M49_U1_nonlinearInst_U6 ( .A1(
        top_AND_M49_U1_nonlinearInst_n50), .A2(
        top_AND_M49_U1_nonlinearInst_n49), .ZN(top_AND_M49_U1_t[0]) );
  AND2_X1 top_AND_M49_U1_nonlinearInst_U5 ( .A1(
        top_AND_M49_U1_nonlinearInst_n48), .A2(
        top_AND_M49_U1_nonlinearInst_n52), .ZN(
        top_AND_M49_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M49_U1_nonlinearInst_U4 ( .A(top_AND_M49_U1_nonlinearInst_n47), .ZN(top_AND_M49_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M49_U1_nonlinearInst_U3 ( .A1(
        top_AND_M49_U1_nonlinearInst_n52), .A2(
        top_AND_M49_U1_nonlinearInst_n48), .ZN(
        top_AND_M49_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M49_U1_nonlinearInst_U2 ( .A1(top_M43), .A2(top_T16), .ZN(
        top_AND_M49_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M49_U1_nonlinearInst_U1 ( .A(Fresh[19]), .ZN(
        top_AND_M49_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M49_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M49_U1_t[0]), .A2(
        top_AND_M49_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M49_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M49_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M49_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M49_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M49_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M49_U1_t_reg[0]) );
  AND2_X1 top_AND_M49_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M49_U1_t[1]), .A2(
        top_AND_M49_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M49_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M49_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M49_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M49_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M49_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M49_U1_t_reg[1]) );
  AND2_X1 top_AND_M49_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M49_U1_t[2]), .A2(
        top_AND_M49_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M49_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M49_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M49_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M49_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M49_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M49_U1_t_reg[2]) );
  AND2_X1 top_AND_M49_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M49_U1_t[3]), .A2(
        top_AND_M49_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M49_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M49_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M49_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M49_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M49_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M49_U1_t_reg[3]) );
  AND2_X1 top_AND_M49_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M49_U1_t[4]), .A2(
        top_AND_M49_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M49_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M49_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M49_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M49_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M49_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M49_U1_t_reg[4]) );
  AND2_X1 top_AND_M49_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M49_U1_t[5]), .A2(
        top_AND_M49_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M49_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M49_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M49_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M49_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M49_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M49_U1_t_reg[5]) );
  AND2_X1 top_AND_M49_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M49_U1_t[6]), .A2(
        top_AND_M49_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M49_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M49_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M49_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M49_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M49_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M49_U1_t_reg[6]) );
  AND2_X1 top_AND_M49_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M49_U1_t[7]), .A2(
        top_AND_M49_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M49_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M49_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M49_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M49_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M49_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M49_U1_t_reg[7]) );
  AND2_X1 top_AND_M49_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_200), .A2(
        top_AND_M49_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M49_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M49_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_310), .A2(top_AND_M49_U1_t_reg[0]), .ZN(
        top_AND_M49_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M49_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_199), .A2(
        top_AND_M49_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M49_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M49_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_310), .A2(top_AND_M49_U1_t_reg[1]), .ZN(
        top_AND_M49_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M49_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_200), .A2(
        top_AND_M49_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M49_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M49_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_309), .A2(top_AND_M49_U1_t_reg[2]), .ZN(
        top_AND_M49_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M49_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_199), .A2(
        top_AND_M49_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M49_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M49_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_309), .A2(top_AND_M49_U1_t_reg[3]), .ZN(
        top_AND_M49_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M49_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M49_U1_OperationInst_q[1]), .A2(
        top_AND_M49_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_333) );
  OR2_X1 top_AND_M49_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M49_U1_OperationInst_q[0]), .A2(
        top_AND_M49_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M49_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M49_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M49_U1_OperationInst_q[3]), .A2(
        top_AND_M49_U1_OperationInst_q[2]), .ZN(
        top_AND_M49_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M49_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_200), .A2(
        top_AND_M49_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M49_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M49_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_310), .A2(top_AND_M49_U1_t_reg[4]), .ZN(
        top_AND_M49_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M49_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_199), .A2(
        top_AND_M49_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M49_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M49_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_310), .A2(top_AND_M49_U1_t_reg[5]), .ZN(
        top_AND_M49_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M49_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_200), .A2(
        top_AND_M49_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M49_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M49_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_309), .A2(top_AND_M49_U1_t_reg[6]), .ZN(
        top_AND_M49_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M49_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_199), .A2(
        top_AND_M49_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M49_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M49_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_309), .A2(top_AND_M49_U1_t_reg[7]), .ZN(
        top_AND_M49_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M49_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M49_U1_OperationInst_q[5]), .A2(
        top_AND_M49_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_334) );
  OR2_X1 top_AND_M49_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M49_U1_OperationInst_q[4]), .A2(
        top_AND_M49_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M49_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M49_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M49_U1_OperationInst_q[7]), .A2(
        top_AND_M49_U1_OperationInst_q[6]), .ZN(
        top_AND_M49_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M50_U1_nonlinearInst_U26 ( .A(top_AND_M50_U1_t[3]), .ZN(
        top_AND_M50_U1_t[7]) );
  OR2_X1 top_AND_M50_U1_nonlinearInst_U25 ( .A1(
        top_AND_M50_U1_nonlinearInst_n64), .A2(
        top_AND_M50_U1_nonlinearInst_n63), .ZN(top_AND_M50_U1_t[3]) );
  INV_X1 top_AND_M50_U1_nonlinearInst_U24 ( .A(
        top_AND_M50_U1_nonlinearInst_n62), .ZN(
        top_AND_M50_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M50_U1_nonlinearInst_U23 ( .A1(
        top_AND_M50_U1_nonlinearInst_n61), .A2(Fresh[20]), .ZN(
        top_AND_M50_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M50_U1_nonlinearInst_U22 ( .A1(Fresh[20]), .A2(
        top_AND_M50_U1_nonlinearInst_n61), .ZN(
        top_AND_M50_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M50_U1_nonlinearInst_U21 ( .A1(top_M38), .A2(top_T9), .ZN(
        top_AND_M50_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M50_U1_nonlinearInst_U20 ( .A(top_AND_M50_U1_t[2]), .ZN(
        top_AND_M50_U1_t[6]) );
  OR2_X1 top_AND_M50_U1_nonlinearInst_U19 ( .A1(
        top_AND_M50_U1_nonlinearInst_n60), .A2(
        top_AND_M50_U1_nonlinearInst_n59), .ZN(top_AND_M50_U1_t[2]) );
  INV_X1 top_AND_M50_U1_nonlinearInst_U18 ( .A(
        top_AND_M50_U1_nonlinearInst_n58), .ZN(
        top_AND_M50_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M50_U1_nonlinearInst_U17 ( .A1(
        top_AND_M50_U1_nonlinearInst_n57), .A2(Fresh[20]), .ZN(
        top_AND_M50_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M50_U1_nonlinearInst_U16 ( .A1(Fresh[20]), .A2(
        top_AND_M50_U1_nonlinearInst_n57), .ZN(
        top_AND_M50_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M50_U1_nonlinearInst_U15 ( .A1(
        top_AND_M50_U1_nonlinearInst_n56), .A2(top_M38), .ZN(
        top_AND_M50_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M50_U1_nonlinearInst_U14 ( .A(top_AND_M50_U1_t[1]), .ZN(
        top_AND_M50_U1_t[5]) );
  OR2_X1 top_AND_M50_U1_nonlinearInst_U13 ( .A1(
        top_AND_M50_U1_nonlinearInst_n55), .A2(
        top_AND_M50_U1_nonlinearInst_n54), .ZN(top_AND_M50_U1_t[1]) );
  AND2_X1 top_AND_M50_U1_nonlinearInst_U12 ( .A1(
        top_AND_M50_U1_nonlinearInst_n53), .A2(
        top_AND_M50_U1_nonlinearInst_n52), .ZN(
        top_AND_M50_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M50_U1_nonlinearInst_U11 ( .A(
        top_AND_M50_U1_nonlinearInst_n51), .ZN(
        top_AND_M50_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M50_U1_nonlinearInst_U10 ( .A1(
        top_AND_M50_U1_nonlinearInst_n52), .A2(
        top_AND_M50_U1_nonlinearInst_n53), .ZN(
        top_AND_M50_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M50_U1_nonlinearInst_U9 ( .A1(top_M38), .A2(
        top_AND_M50_U1_nonlinearInst_n56), .ZN(
        top_AND_M50_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M50_U1_nonlinearInst_U8 ( .A(top_T9), .ZN(
        top_AND_M50_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M50_U1_nonlinearInst_U7 ( .A(top_AND_M50_U1_t[0]), .ZN(
        top_AND_M50_U1_t[4]) );
  OR2_X1 top_AND_M50_U1_nonlinearInst_U6 ( .A1(
        top_AND_M50_U1_nonlinearInst_n50), .A2(
        top_AND_M50_U1_nonlinearInst_n49), .ZN(top_AND_M50_U1_t[0]) );
  AND2_X1 top_AND_M50_U1_nonlinearInst_U5 ( .A1(
        top_AND_M50_U1_nonlinearInst_n48), .A2(
        top_AND_M50_U1_nonlinearInst_n52), .ZN(
        top_AND_M50_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M50_U1_nonlinearInst_U4 ( .A(top_AND_M50_U1_nonlinearInst_n47), .ZN(top_AND_M50_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M50_U1_nonlinearInst_U3 ( .A1(
        top_AND_M50_U1_nonlinearInst_n52), .A2(
        top_AND_M50_U1_nonlinearInst_n48), .ZN(
        top_AND_M50_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M50_U1_nonlinearInst_U2 ( .A1(top_M38), .A2(top_T9), .ZN(
        top_AND_M50_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M50_U1_nonlinearInst_U1 ( .A(Fresh[20]), .ZN(
        top_AND_M50_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M50_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M50_U1_t[0]), .A2(
        top_AND_M50_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M50_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M50_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M50_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M50_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M50_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M50_U1_t_reg[0]) );
  AND2_X1 top_AND_M50_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M50_U1_t[1]), .A2(
        top_AND_M50_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M50_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M50_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M50_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M50_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M50_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M50_U1_t_reg[1]) );
  AND2_X1 top_AND_M50_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M50_U1_t[2]), .A2(
        top_AND_M50_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M50_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M50_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M50_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M50_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M50_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M50_U1_t_reg[2]) );
  AND2_X1 top_AND_M50_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M50_U1_t[3]), .A2(
        top_AND_M50_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M50_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M50_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M50_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M50_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M50_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M50_U1_t_reg[3]) );
  AND2_X1 top_AND_M50_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M50_U1_t[4]), .A2(
        top_AND_M50_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M50_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M50_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M50_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M50_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M50_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M50_U1_t_reg[4]) );
  AND2_X1 top_AND_M50_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M50_U1_t[5]), .A2(
        top_AND_M50_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M50_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M50_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M50_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M50_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M50_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M50_U1_t_reg[5]) );
  AND2_X1 top_AND_M50_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M50_U1_t[6]), .A2(
        top_AND_M50_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M50_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M50_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M50_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M50_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M50_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M50_U1_t_reg[6]) );
  AND2_X1 top_AND_M50_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M50_U1_t[7]), .A2(
        top_AND_M50_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M50_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M50_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M50_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M50_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M50_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M50_U1_t_reg[7]) );
  AND2_X1 top_AND_M50_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_194), .A2(
        top_AND_M50_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M50_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M50_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_300), .A2(top_AND_M50_U1_t_reg[0]), .ZN(
        top_AND_M50_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M50_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_193), .A2(
        top_AND_M50_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M50_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M50_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_300), .A2(top_AND_M50_U1_t_reg[1]), .ZN(
        top_AND_M50_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M50_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_194), .A2(
        top_AND_M50_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M50_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M50_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_299), .A2(top_AND_M50_U1_t_reg[2]), .ZN(
        top_AND_M50_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M50_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_193), .A2(
        top_AND_M50_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M50_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M50_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_299), .A2(top_AND_M50_U1_t_reg[3]), .ZN(
        top_AND_M50_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M50_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M50_U1_OperationInst_q[1]), .A2(
        top_AND_M50_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_317) );
  OR2_X1 top_AND_M50_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M50_U1_OperationInst_q[0]), .A2(
        top_AND_M50_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M50_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M50_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M50_U1_OperationInst_q[3]), .A2(
        top_AND_M50_U1_OperationInst_q[2]), .ZN(
        top_AND_M50_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M50_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_194), .A2(
        top_AND_M50_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M50_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M50_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_300), .A2(top_AND_M50_U1_t_reg[4]), .ZN(
        top_AND_M50_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M50_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_193), .A2(
        top_AND_M50_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M50_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M50_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_300), .A2(top_AND_M50_U1_t_reg[5]), .ZN(
        top_AND_M50_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M50_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_194), .A2(
        top_AND_M50_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M50_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M50_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_299), .A2(top_AND_M50_U1_t_reg[6]), .ZN(
        top_AND_M50_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M50_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_193), .A2(
        top_AND_M50_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M50_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M50_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_299), .A2(top_AND_M50_U1_t_reg[7]), .ZN(
        top_AND_M50_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M50_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M50_U1_OperationInst_q[5]), .A2(
        top_AND_M50_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_318) );
  OR2_X1 top_AND_M50_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M50_U1_OperationInst_q[4]), .A2(
        top_AND_M50_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M50_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M50_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M50_U1_OperationInst_q[7]), .A2(
        top_AND_M50_U1_OperationInst_q[6]), .ZN(
        top_AND_M50_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M51_U1_nonlinearInst_U26 ( .A(top_AND_M51_U1_t[3]), .ZN(
        top_AND_M51_U1_t[7]) );
  OR2_X1 top_AND_M51_U1_nonlinearInst_U25 ( .A1(
        top_AND_M51_U1_nonlinearInst_n64), .A2(
        top_AND_M51_U1_nonlinearInst_n63), .ZN(top_AND_M51_U1_t[3]) );
  INV_X1 top_AND_M51_U1_nonlinearInst_U24 ( .A(
        top_AND_M51_U1_nonlinearInst_n62), .ZN(
        top_AND_M51_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M51_U1_nonlinearInst_U23 ( .A1(
        top_AND_M51_U1_nonlinearInst_n61), .A2(Fresh[21]), .ZN(
        top_AND_M51_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M51_U1_nonlinearInst_U22 ( .A1(Fresh[21]), .A2(
        top_AND_M51_U1_nonlinearInst_n61), .ZN(
        top_AND_M51_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M51_U1_nonlinearInst_U21 ( .A1(top_M37), .A2(top_T17), .ZN(
        top_AND_M51_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M51_U1_nonlinearInst_U20 ( .A(top_AND_M51_U1_t[2]), .ZN(
        top_AND_M51_U1_t[6]) );
  OR2_X1 top_AND_M51_U1_nonlinearInst_U19 ( .A1(
        top_AND_M51_U1_nonlinearInst_n60), .A2(
        top_AND_M51_U1_nonlinearInst_n59), .ZN(top_AND_M51_U1_t[2]) );
  INV_X1 top_AND_M51_U1_nonlinearInst_U18 ( .A(
        top_AND_M51_U1_nonlinearInst_n58), .ZN(
        top_AND_M51_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M51_U1_nonlinearInst_U17 ( .A1(
        top_AND_M51_U1_nonlinearInst_n57), .A2(Fresh[21]), .ZN(
        top_AND_M51_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M51_U1_nonlinearInst_U16 ( .A1(Fresh[21]), .A2(
        top_AND_M51_U1_nonlinearInst_n57), .ZN(
        top_AND_M51_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M51_U1_nonlinearInst_U15 ( .A1(
        top_AND_M51_U1_nonlinearInst_n56), .A2(top_M37), .ZN(
        top_AND_M51_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M51_U1_nonlinearInst_U14 ( .A(top_AND_M51_U1_t[1]), .ZN(
        top_AND_M51_U1_t[5]) );
  OR2_X1 top_AND_M51_U1_nonlinearInst_U13 ( .A1(
        top_AND_M51_U1_nonlinearInst_n55), .A2(
        top_AND_M51_U1_nonlinearInst_n54), .ZN(top_AND_M51_U1_t[1]) );
  AND2_X1 top_AND_M51_U1_nonlinearInst_U12 ( .A1(
        top_AND_M51_U1_nonlinearInst_n53), .A2(
        top_AND_M51_U1_nonlinearInst_n52), .ZN(
        top_AND_M51_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M51_U1_nonlinearInst_U11 ( .A(
        top_AND_M51_U1_nonlinearInst_n51), .ZN(
        top_AND_M51_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M51_U1_nonlinearInst_U10 ( .A1(
        top_AND_M51_U1_nonlinearInst_n52), .A2(
        top_AND_M51_U1_nonlinearInst_n53), .ZN(
        top_AND_M51_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M51_U1_nonlinearInst_U9 ( .A1(top_M37), .A2(
        top_AND_M51_U1_nonlinearInst_n56), .ZN(
        top_AND_M51_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M51_U1_nonlinearInst_U8 ( .A(top_T17), .ZN(
        top_AND_M51_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M51_U1_nonlinearInst_U7 ( .A(top_AND_M51_U1_t[0]), .ZN(
        top_AND_M51_U1_t[4]) );
  OR2_X1 top_AND_M51_U1_nonlinearInst_U6 ( .A1(
        top_AND_M51_U1_nonlinearInst_n50), .A2(
        top_AND_M51_U1_nonlinearInst_n49), .ZN(top_AND_M51_U1_t[0]) );
  AND2_X1 top_AND_M51_U1_nonlinearInst_U5 ( .A1(
        top_AND_M51_U1_nonlinearInst_n48), .A2(
        top_AND_M51_U1_nonlinearInst_n52), .ZN(
        top_AND_M51_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M51_U1_nonlinearInst_U4 ( .A(top_AND_M51_U1_nonlinearInst_n47), .ZN(top_AND_M51_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M51_U1_nonlinearInst_U3 ( .A1(
        top_AND_M51_U1_nonlinearInst_n52), .A2(
        top_AND_M51_U1_nonlinearInst_n48), .ZN(
        top_AND_M51_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M51_U1_nonlinearInst_U2 ( .A1(top_M37), .A2(top_T17), .ZN(
        top_AND_M51_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M51_U1_nonlinearInst_U1 ( .A(Fresh[21]), .ZN(
        top_AND_M51_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M51_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M51_U1_t[0]), .A2(
        top_AND_M51_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M51_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M51_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M51_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M51_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M51_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M51_U1_t_reg[0]) );
  AND2_X1 top_AND_M51_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M51_U1_t[1]), .A2(
        top_AND_M51_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M51_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M51_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M51_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M51_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M51_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M51_U1_t_reg[1]) );
  AND2_X1 top_AND_M51_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M51_U1_t[2]), .A2(
        top_AND_M51_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M51_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M51_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M51_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M51_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M51_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M51_U1_t_reg[2]) );
  AND2_X1 top_AND_M51_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M51_U1_t[3]), .A2(
        top_AND_M51_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M51_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M51_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M51_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M51_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M51_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M51_U1_t_reg[3]) );
  AND2_X1 top_AND_M51_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M51_U1_t[4]), .A2(
        top_AND_M51_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M51_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M51_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M51_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M51_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M51_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M51_U1_t_reg[4]) );
  AND2_X1 top_AND_M51_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M51_U1_t[5]), .A2(
        top_AND_M51_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M51_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M51_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M51_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M51_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M51_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M51_U1_t_reg[5]) );
  AND2_X1 top_AND_M51_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M51_U1_t[6]), .A2(
        top_AND_M51_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M51_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M51_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M51_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M51_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M51_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M51_U1_t_reg[6]) );
  AND2_X1 top_AND_M51_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M51_U1_t[7]), .A2(
        top_AND_M51_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M51_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M51_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M51_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M51_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M51_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M51_U1_t_reg[7]) );
  AND2_X1 top_AND_M51_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_214), .A2(
        top_AND_M51_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M51_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M51_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_298), .A2(top_AND_M51_U1_t_reg[0]), .ZN(
        top_AND_M51_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M51_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_213), .A2(
        top_AND_M51_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M51_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M51_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_298), .A2(top_AND_M51_U1_t_reg[1]), .ZN(
        top_AND_M51_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M51_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_214), .A2(
        top_AND_M51_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M51_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M51_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_297), .A2(top_AND_M51_U1_t_reg[2]), .ZN(
        top_AND_M51_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M51_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_213), .A2(
        top_AND_M51_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M51_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M51_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_297), .A2(top_AND_M51_U1_t_reg[3]), .ZN(
        top_AND_M51_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M51_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M51_U1_OperationInst_q[1]), .A2(
        top_AND_M51_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_319) );
  OR2_X1 top_AND_M51_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M51_U1_OperationInst_q[0]), .A2(
        top_AND_M51_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M51_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M51_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M51_U1_OperationInst_q[3]), .A2(
        top_AND_M51_U1_OperationInst_q[2]), .ZN(
        top_AND_M51_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M51_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_214), .A2(
        top_AND_M51_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M51_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M51_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_298), .A2(top_AND_M51_U1_t_reg[4]), .ZN(
        top_AND_M51_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M51_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_213), .A2(
        top_AND_M51_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M51_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M51_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_298), .A2(top_AND_M51_U1_t_reg[5]), .ZN(
        top_AND_M51_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M51_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_214), .A2(
        top_AND_M51_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M51_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M51_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_297), .A2(top_AND_M51_U1_t_reg[6]), .ZN(
        top_AND_M51_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M51_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_213), .A2(
        top_AND_M51_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M51_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M51_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_297), .A2(top_AND_M51_U1_t_reg[7]), .ZN(
        top_AND_M51_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M51_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M51_U1_OperationInst_q[5]), .A2(
        top_AND_M51_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_320) );
  OR2_X1 top_AND_M51_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M51_U1_OperationInst_q[4]), .A2(
        top_AND_M51_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M51_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M51_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M51_U1_OperationInst_q[7]), .A2(
        top_AND_M51_U1_OperationInst_q[6]), .ZN(
        top_AND_M51_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M52_U1_nonlinearInst_U26 ( .A(top_AND_M52_U1_t[3]), .ZN(
        top_AND_M52_U1_t[7]) );
  OR2_X1 top_AND_M52_U1_nonlinearInst_U25 ( .A1(
        top_AND_M52_U1_nonlinearInst_n64), .A2(
        top_AND_M52_U1_nonlinearInst_n63), .ZN(top_AND_M52_U1_t[3]) );
  INV_X1 top_AND_M52_U1_nonlinearInst_U24 ( .A(
        top_AND_M52_U1_nonlinearInst_n62), .ZN(
        top_AND_M52_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M52_U1_nonlinearInst_U23 ( .A1(
        top_AND_M52_U1_nonlinearInst_n61), .A2(Fresh[22]), .ZN(
        top_AND_M52_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M52_U1_nonlinearInst_U22 ( .A1(Fresh[22]), .A2(
        top_AND_M52_U1_nonlinearInst_n61), .ZN(
        top_AND_M52_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M52_U1_nonlinearInst_U21 ( .A1(top_M42), .A2(top_T15), .ZN(
        top_AND_M52_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M52_U1_nonlinearInst_U20 ( .A(top_AND_M52_U1_t[2]), .ZN(
        top_AND_M52_U1_t[6]) );
  OR2_X1 top_AND_M52_U1_nonlinearInst_U19 ( .A1(
        top_AND_M52_U1_nonlinearInst_n60), .A2(
        top_AND_M52_U1_nonlinearInst_n59), .ZN(top_AND_M52_U1_t[2]) );
  INV_X1 top_AND_M52_U1_nonlinearInst_U18 ( .A(
        top_AND_M52_U1_nonlinearInst_n58), .ZN(
        top_AND_M52_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M52_U1_nonlinearInst_U17 ( .A1(
        top_AND_M52_U1_nonlinearInst_n57), .A2(Fresh[22]), .ZN(
        top_AND_M52_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M52_U1_nonlinearInst_U16 ( .A1(Fresh[22]), .A2(
        top_AND_M52_U1_nonlinearInst_n57), .ZN(
        top_AND_M52_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M52_U1_nonlinearInst_U15 ( .A1(
        top_AND_M52_U1_nonlinearInst_n56), .A2(top_M42), .ZN(
        top_AND_M52_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M52_U1_nonlinearInst_U14 ( .A(top_AND_M52_U1_t[1]), .ZN(
        top_AND_M52_U1_t[5]) );
  OR2_X1 top_AND_M52_U1_nonlinearInst_U13 ( .A1(
        top_AND_M52_U1_nonlinearInst_n55), .A2(
        top_AND_M52_U1_nonlinearInst_n54), .ZN(top_AND_M52_U1_t[1]) );
  AND2_X1 top_AND_M52_U1_nonlinearInst_U12 ( .A1(
        top_AND_M52_U1_nonlinearInst_n53), .A2(
        top_AND_M52_U1_nonlinearInst_n52), .ZN(
        top_AND_M52_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M52_U1_nonlinearInst_U11 ( .A(
        top_AND_M52_U1_nonlinearInst_n51), .ZN(
        top_AND_M52_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M52_U1_nonlinearInst_U10 ( .A1(
        top_AND_M52_U1_nonlinearInst_n52), .A2(
        top_AND_M52_U1_nonlinearInst_n53), .ZN(
        top_AND_M52_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M52_U1_nonlinearInst_U9 ( .A1(top_M42), .A2(
        top_AND_M52_U1_nonlinearInst_n56), .ZN(
        top_AND_M52_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M52_U1_nonlinearInst_U8 ( .A(top_T15), .ZN(
        top_AND_M52_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M52_U1_nonlinearInst_U7 ( .A(top_AND_M52_U1_t[0]), .ZN(
        top_AND_M52_U1_t[4]) );
  OR2_X1 top_AND_M52_U1_nonlinearInst_U6 ( .A1(
        top_AND_M52_U1_nonlinearInst_n50), .A2(
        top_AND_M52_U1_nonlinearInst_n49), .ZN(top_AND_M52_U1_t[0]) );
  AND2_X1 top_AND_M52_U1_nonlinearInst_U5 ( .A1(
        top_AND_M52_U1_nonlinearInst_n48), .A2(
        top_AND_M52_U1_nonlinearInst_n52), .ZN(
        top_AND_M52_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M52_U1_nonlinearInst_U4 ( .A(top_AND_M52_U1_nonlinearInst_n47), .ZN(top_AND_M52_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M52_U1_nonlinearInst_U3 ( .A1(
        top_AND_M52_U1_nonlinearInst_n52), .A2(
        top_AND_M52_U1_nonlinearInst_n48), .ZN(
        top_AND_M52_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M52_U1_nonlinearInst_U2 ( .A1(top_M42), .A2(top_T15), .ZN(
        top_AND_M52_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M52_U1_nonlinearInst_U1 ( .A(Fresh[22]), .ZN(
        top_AND_M52_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M52_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M52_U1_t[0]), .A2(
        top_AND_M52_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M52_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M52_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M52_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M52_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M52_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M52_U1_t_reg[0]) );
  AND2_X1 top_AND_M52_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M52_U1_t[1]), .A2(
        top_AND_M52_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M52_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M52_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M52_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M52_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M52_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M52_U1_t_reg[1]) );
  AND2_X1 top_AND_M52_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M52_U1_t[2]), .A2(
        top_AND_M52_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M52_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M52_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M52_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M52_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M52_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M52_U1_t_reg[2]) );
  AND2_X1 top_AND_M52_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M52_U1_t[3]), .A2(
        top_AND_M52_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M52_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M52_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M52_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M52_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M52_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M52_U1_t_reg[3]) );
  AND2_X1 top_AND_M52_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M52_U1_t[4]), .A2(
        top_AND_M52_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M52_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M52_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M52_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M52_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M52_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M52_U1_t_reg[4]) );
  AND2_X1 top_AND_M52_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M52_U1_t[5]), .A2(
        top_AND_M52_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M52_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M52_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M52_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M52_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M52_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M52_U1_t_reg[5]) );
  AND2_X1 top_AND_M52_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M52_U1_t[6]), .A2(
        top_AND_M52_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M52_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M52_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M52_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M52_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M52_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M52_U1_t_reg[6]) );
  AND2_X1 top_AND_M52_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M52_U1_t[7]), .A2(
        top_AND_M52_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M52_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M52_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M52_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M52_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M52_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M52_U1_t_reg[7]) );
  AND2_X1 top_AND_M52_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_198), .A2(
        top_AND_M52_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M52_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M52_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_308), .A2(top_AND_M52_U1_t_reg[0]), .ZN(
        top_AND_M52_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M52_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_197), .A2(
        top_AND_M52_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M52_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M52_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_308), .A2(top_AND_M52_U1_t_reg[1]), .ZN(
        top_AND_M52_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M52_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_198), .A2(
        top_AND_M52_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M52_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M52_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_307), .A2(top_AND_M52_U1_t_reg[2]), .ZN(
        top_AND_M52_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M52_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_197), .A2(
        top_AND_M52_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M52_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M52_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_307), .A2(top_AND_M52_U1_t_reg[3]), .ZN(
        top_AND_M52_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M52_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M52_U1_OperationInst_q[1]), .A2(
        top_AND_M52_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_335) );
  OR2_X1 top_AND_M52_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M52_U1_OperationInst_q[0]), .A2(
        top_AND_M52_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M52_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M52_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M52_U1_OperationInst_q[3]), .A2(
        top_AND_M52_U1_OperationInst_q[2]), .ZN(
        top_AND_M52_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M52_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_198), .A2(
        top_AND_M52_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M52_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M52_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_308), .A2(top_AND_M52_U1_t_reg[4]), .ZN(
        top_AND_M52_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M52_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_197), .A2(
        top_AND_M52_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M52_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M52_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_308), .A2(top_AND_M52_U1_t_reg[5]), .ZN(
        top_AND_M52_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M52_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_198), .A2(
        top_AND_M52_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M52_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M52_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_307), .A2(top_AND_M52_U1_t_reg[6]), .ZN(
        top_AND_M52_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M52_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_197), .A2(
        top_AND_M52_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M52_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M52_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_307), .A2(top_AND_M52_U1_t_reg[7]), .ZN(
        top_AND_M52_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M52_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M52_U1_OperationInst_q[5]), .A2(
        top_AND_M52_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_336) );
  OR2_X1 top_AND_M52_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M52_U1_OperationInst_q[4]), .A2(
        top_AND_M52_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M52_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M52_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M52_U1_OperationInst_q[7]), .A2(
        top_AND_M52_U1_OperationInst_q[6]), .ZN(
        top_AND_M52_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M53_U1_nonlinearInst_U26 ( .A(top_AND_M53_U1_t[3]), .ZN(
        top_AND_M53_U1_t[7]) );
  OR2_X1 top_AND_M53_U1_nonlinearInst_U25 ( .A1(
        top_AND_M53_U1_nonlinearInst_n64), .A2(
        top_AND_M53_U1_nonlinearInst_n63), .ZN(top_AND_M53_U1_t[3]) );
  INV_X1 top_AND_M53_U1_nonlinearInst_U24 ( .A(
        top_AND_M53_U1_nonlinearInst_n62), .ZN(
        top_AND_M53_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M53_U1_nonlinearInst_U23 ( .A1(
        top_AND_M53_U1_nonlinearInst_n61), .A2(Fresh[23]), .ZN(
        top_AND_M53_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M53_U1_nonlinearInst_U22 ( .A1(Fresh[23]), .A2(
        top_AND_M53_U1_nonlinearInst_n61), .ZN(
        top_AND_M53_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M53_U1_nonlinearInst_U21 ( .A1(top_M45), .A2(top_T27), .ZN(
        top_AND_M53_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M53_U1_nonlinearInst_U20 ( .A(top_AND_M53_U1_t[2]), .ZN(
        top_AND_M53_U1_t[6]) );
  OR2_X1 top_AND_M53_U1_nonlinearInst_U19 ( .A1(
        top_AND_M53_U1_nonlinearInst_n60), .A2(
        top_AND_M53_U1_nonlinearInst_n59), .ZN(top_AND_M53_U1_t[2]) );
  INV_X1 top_AND_M53_U1_nonlinearInst_U18 ( .A(
        top_AND_M53_U1_nonlinearInst_n58), .ZN(
        top_AND_M53_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M53_U1_nonlinearInst_U17 ( .A1(
        top_AND_M53_U1_nonlinearInst_n57), .A2(Fresh[23]), .ZN(
        top_AND_M53_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M53_U1_nonlinearInst_U16 ( .A1(Fresh[23]), .A2(
        top_AND_M53_U1_nonlinearInst_n57), .ZN(
        top_AND_M53_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M53_U1_nonlinearInst_U15 ( .A1(
        top_AND_M53_U1_nonlinearInst_n56), .A2(top_M45), .ZN(
        top_AND_M53_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M53_U1_nonlinearInst_U14 ( .A(top_AND_M53_U1_t[1]), .ZN(
        top_AND_M53_U1_t[5]) );
  OR2_X1 top_AND_M53_U1_nonlinearInst_U13 ( .A1(
        top_AND_M53_U1_nonlinearInst_n55), .A2(
        top_AND_M53_U1_nonlinearInst_n54), .ZN(top_AND_M53_U1_t[1]) );
  AND2_X1 top_AND_M53_U1_nonlinearInst_U12 ( .A1(
        top_AND_M53_U1_nonlinearInst_n53), .A2(
        top_AND_M53_U1_nonlinearInst_n52), .ZN(
        top_AND_M53_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M53_U1_nonlinearInst_U11 ( .A(
        top_AND_M53_U1_nonlinearInst_n51), .ZN(
        top_AND_M53_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M53_U1_nonlinearInst_U10 ( .A1(
        top_AND_M53_U1_nonlinearInst_n52), .A2(
        top_AND_M53_U1_nonlinearInst_n53), .ZN(
        top_AND_M53_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M53_U1_nonlinearInst_U9 ( .A1(top_M45), .A2(
        top_AND_M53_U1_nonlinearInst_n56), .ZN(
        top_AND_M53_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M53_U1_nonlinearInst_U8 ( .A(top_T27), .ZN(
        top_AND_M53_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M53_U1_nonlinearInst_U7 ( .A(top_AND_M53_U1_t[0]), .ZN(
        top_AND_M53_U1_t[4]) );
  OR2_X1 top_AND_M53_U1_nonlinearInst_U6 ( .A1(
        top_AND_M53_U1_nonlinearInst_n50), .A2(
        top_AND_M53_U1_nonlinearInst_n49), .ZN(top_AND_M53_U1_t[0]) );
  AND2_X1 top_AND_M53_U1_nonlinearInst_U5 ( .A1(
        top_AND_M53_U1_nonlinearInst_n48), .A2(
        top_AND_M53_U1_nonlinearInst_n52), .ZN(
        top_AND_M53_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M53_U1_nonlinearInst_U4 ( .A(top_AND_M53_U1_nonlinearInst_n47), .ZN(top_AND_M53_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M53_U1_nonlinearInst_U3 ( .A1(
        top_AND_M53_U1_nonlinearInst_n52), .A2(
        top_AND_M53_U1_nonlinearInst_n48), .ZN(
        top_AND_M53_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M53_U1_nonlinearInst_U2 ( .A1(top_M45), .A2(top_T27), .ZN(
        top_AND_M53_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M53_U1_nonlinearInst_U1 ( .A(Fresh[23]), .ZN(
        top_AND_M53_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M53_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M53_U1_t[0]), .A2(
        top_AND_M53_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M53_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M53_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M53_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M53_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M53_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M53_U1_t_reg[0]) );
  AND2_X1 top_AND_M53_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M53_U1_t[1]), .A2(
        top_AND_M53_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M53_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M53_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M53_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M53_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M53_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M53_U1_t_reg[1]) );
  AND2_X1 top_AND_M53_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M53_U1_t[2]), .A2(
        top_AND_M53_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M53_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M53_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M53_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M53_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M53_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M53_U1_t_reg[2]) );
  AND2_X1 top_AND_M53_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M53_U1_t[3]), .A2(
        top_AND_M53_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M53_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M53_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M53_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M53_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M53_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M53_U1_t_reg[3]) );
  AND2_X1 top_AND_M53_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M53_U1_t[4]), .A2(
        top_AND_M53_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M53_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M53_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M53_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M53_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M53_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M53_U1_t_reg[4]) );
  AND2_X1 top_AND_M53_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M53_U1_t[5]), .A2(
        top_AND_M53_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M53_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M53_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M53_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M53_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M53_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M53_U1_t_reg[5]) );
  AND2_X1 top_AND_M53_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M53_U1_t[6]), .A2(
        top_AND_M53_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M53_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M53_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M53_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M53_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M53_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M53_U1_t_reg[6]) );
  AND2_X1 top_AND_M53_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M53_U1_t[7]), .A2(
        top_AND_M53_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M53_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M53_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M53_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M53_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M53_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M53_U1_t_reg[7]) );
  AND2_X1 top_AND_M53_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_206), .A2(
        top_AND_M53_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M53_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M53_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_330), .A2(top_AND_M53_U1_t_reg[0]), .ZN(
        top_AND_M53_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M53_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_205), .A2(
        top_AND_M53_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M53_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M53_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_330), .A2(top_AND_M53_U1_t_reg[1]), .ZN(
        top_AND_M53_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M53_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_206), .A2(
        top_AND_M53_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M53_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M53_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_329), .A2(top_AND_M53_U1_t_reg[2]), .ZN(
        top_AND_M53_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M53_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_205), .A2(
        top_AND_M53_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M53_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M53_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_329), .A2(top_AND_M53_U1_t_reg[3]), .ZN(
        top_AND_M53_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M53_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M53_U1_OperationInst_q[1]), .A2(
        top_AND_M53_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_353) );
  OR2_X1 top_AND_M53_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M53_U1_OperationInst_q[0]), .A2(
        top_AND_M53_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M53_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M53_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M53_U1_OperationInst_q[3]), .A2(
        top_AND_M53_U1_OperationInst_q[2]), .ZN(
        top_AND_M53_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M53_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_206), .A2(
        top_AND_M53_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M53_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M53_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_330), .A2(top_AND_M53_U1_t_reg[4]), .ZN(
        top_AND_M53_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M53_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_205), .A2(
        top_AND_M53_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M53_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M53_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_330), .A2(top_AND_M53_U1_t_reg[5]), .ZN(
        top_AND_M53_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M53_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_206), .A2(
        top_AND_M53_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M53_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M53_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_329), .A2(top_AND_M53_U1_t_reg[6]), .ZN(
        top_AND_M53_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M53_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_205), .A2(
        top_AND_M53_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M53_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M53_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_329), .A2(top_AND_M53_U1_t_reg[7]), .ZN(
        top_AND_M53_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M53_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M53_U1_OperationInst_q[5]), .A2(
        top_AND_M53_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_354) );
  OR2_X1 top_AND_M53_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M53_U1_OperationInst_q[4]), .A2(
        top_AND_M53_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M53_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M53_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M53_U1_OperationInst_q[7]), .A2(
        top_AND_M53_U1_OperationInst_q[6]), .ZN(
        top_AND_M53_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M54_U1_nonlinearInst_U26 ( .A(top_AND_M54_U1_t[3]), .ZN(
        top_AND_M54_U1_t[7]) );
  OR2_X1 top_AND_M54_U1_nonlinearInst_U25 ( .A1(
        top_AND_M54_U1_nonlinearInst_n64), .A2(
        top_AND_M54_U1_nonlinearInst_n63), .ZN(top_AND_M54_U1_t[3]) );
  INV_X1 top_AND_M54_U1_nonlinearInst_U24 ( .A(
        top_AND_M54_U1_nonlinearInst_n62), .ZN(
        top_AND_M54_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M54_U1_nonlinearInst_U23 ( .A1(
        top_AND_M54_U1_nonlinearInst_n61), .A2(Fresh[24]), .ZN(
        top_AND_M54_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M54_U1_nonlinearInst_U22 ( .A1(Fresh[24]), .A2(
        top_AND_M54_U1_nonlinearInst_n61), .ZN(
        top_AND_M54_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M54_U1_nonlinearInst_U21 ( .A1(top_M41), .A2(top_T10), .ZN(
        top_AND_M54_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M54_U1_nonlinearInst_U20 ( .A(top_AND_M54_U1_t[2]), .ZN(
        top_AND_M54_U1_t[6]) );
  OR2_X1 top_AND_M54_U1_nonlinearInst_U19 ( .A1(
        top_AND_M54_U1_nonlinearInst_n60), .A2(
        top_AND_M54_U1_nonlinearInst_n59), .ZN(top_AND_M54_U1_t[2]) );
  INV_X1 top_AND_M54_U1_nonlinearInst_U18 ( .A(
        top_AND_M54_U1_nonlinearInst_n58), .ZN(
        top_AND_M54_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M54_U1_nonlinearInst_U17 ( .A1(
        top_AND_M54_U1_nonlinearInst_n57), .A2(Fresh[24]), .ZN(
        top_AND_M54_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M54_U1_nonlinearInst_U16 ( .A1(Fresh[24]), .A2(
        top_AND_M54_U1_nonlinearInst_n57), .ZN(
        top_AND_M54_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M54_U1_nonlinearInst_U15 ( .A1(
        top_AND_M54_U1_nonlinearInst_n56), .A2(top_M41), .ZN(
        top_AND_M54_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M54_U1_nonlinearInst_U14 ( .A(top_AND_M54_U1_t[1]), .ZN(
        top_AND_M54_U1_t[5]) );
  OR2_X1 top_AND_M54_U1_nonlinearInst_U13 ( .A1(
        top_AND_M54_U1_nonlinearInst_n55), .A2(
        top_AND_M54_U1_nonlinearInst_n54), .ZN(top_AND_M54_U1_t[1]) );
  AND2_X1 top_AND_M54_U1_nonlinearInst_U12 ( .A1(
        top_AND_M54_U1_nonlinearInst_n53), .A2(
        top_AND_M54_U1_nonlinearInst_n52), .ZN(
        top_AND_M54_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M54_U1_nonlinearInst_U11 ( .A(
        top_AND_M54_U1_nonlinearInst_n51), .ZN(
        top_AND_M54_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M54_U1_nonlinearInst_U10 ( .A1(
        top_AND_M54_U1_nonlinearInst_n52), .A2(
        top_AND_M54_U1_nonlinearInst_n53), .ZN(
        top_AND_M54_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M54_U1_nonlinearInst_U9 ( .A1(top_M41), .A2(
        top_AND_M54_U1_nonlinearInst_n56), .ZN(
        top_AND_M54_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M54_U1_nonlinearInst_U8 ( .A(top_T10), .ZN(
        top_AND_M54_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M54_U1_nonlinearInst_U7 ( .A(top_AND_M54_U1_t[0]), .ZN(
        top_AND_M54_U1_t[4]) );
  OR2_X1 top_AND_M54_U1_nonlinearInst_U6 ( .A1(
        top_AND_M54_U1_nonlinearInst_n50), .A2(
        top_AND_M54_U1_nonlinearInst_n49), .ZN(top_AND_M54_U1_t[0]) );
  AND2_X1 top_AND_M54_U1_nonlinearInst_U5 ( .A1(
        top_AND_M54_U1_nonlinearInst_n48), .A2(
        top_AND_M54_U1_nonlinearInst_n52), .ZN(
        top_AND_M54_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M54_U1_nonlinearInst_U4 ( .A(top_AND_M54_U1_nonlinearInst_n47), .ZN(top_AND_M54_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M54_U1_nonlinearInst_U3 ( .A1(
        top_AND_M54_U1_nonlinearInst_n52), .A2(
        top_AND_M54_U1_nonlinearInst_n48), .ZN(
        top_AND_M54_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M54_U1_nonlinearInst_U2 ( .A1(top_M41), .A2(top_T10), .ZN(
        top_AND_M54_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M54_U1_nonlinearInst_U1 ( .A(Fresh[24]), .ZN(
        top_AND_M54_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M54_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M54_U1_t[0]), .A2(
        top_AND_M54_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M54_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M54_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M54_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M54_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M54_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M54_U1_t_reg[0]) );
  AND2_X1 top_AND_M54_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M54_U1_t[1]), .A2(
        top_AND_M54_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M54_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M54_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M54_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M54_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M54_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M54_U1_t_reg[1]) );
  AND2_X1 top_AND_M54_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M54_U1_t[2]), .A2(
        top_AND_M54_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M54_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M54_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M54_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M54_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M54_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M54_U1_t_reg[2]) );
  AND2_X1 top_AND_M54_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M54_U1_t[3]), .A2(
        top_AND_M54_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M54_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M54_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M54_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M54_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M54_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M54_U1_t_reg[3]) );
  AND2_X1 top_AND_M54_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M54_U1_t[4]), .A2(
        top_AND_M54_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M54_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M54_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M54_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M54_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M54_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M54_U1_t_reg[4]) );
  AND2_X1 top_AND_M54_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M54_U1_t[5]), .A2(
        top_AND_M54_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M54_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M54_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M54_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M54_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M54_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M54_U1_t_reg[5]) );
  AND2_X1 top_AND_M54_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M54_U1_t[6]), .A2(
        top_AND_M54_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M54_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M54_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M54_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M54_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M54_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M54_U1_t_reg[6]) );
  AND2_X1 top_AND_M54_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M54_U1_t[7]), .A2(
        top_AND_M54_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M54_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M54_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M54_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M54_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M54_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M54_U1_t_reg[7]) );
  AND2_X1 top_AND_M54_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_210), .A2(
        top_AND_M54_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M54_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M54_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_306), .A2(top_AND_M54_U1_t_reg[0]), .ZN(
        top_AND_M54_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M54_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_209), .A2(
        top_AND_M54_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M54_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M54_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_306), .A2(top_AND_M54_U1_t_reg[1]), .ZN(
        top_AND_M54_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M54_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_210), .A2(
        top_AND_M54_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M54_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M54_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_305), .A2(top_AND_M54_U1_t_reg[2]), .ZN(
        top_AND_M54_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M54_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_209), .A2(
        top_AND_M54_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M54_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M54_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_305), .A2(top_AND_M54_U1_t_reg[3]), .ZN(
        top_AND_M54_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M54_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M54_U1_OperationInst_q[1]), .A2(
        top_AND_M54_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_337) );
  OR2_X1 top_AND_M54_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M54_U1_OperationInst_q[0]), .A2(
        top_AND_M54_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M54_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M54_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M54_U1_OperationInst_q[3]), .A2(
        top_AND_M54_U1_OperationInst_q[2]), .ZN(
        top_AND_M54_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M54_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_210), .A2(
        top_AND_M54_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M54_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M54_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_306), .A2(top_AND_M54_U1_t_reg[4]), .ZN(
        top_AND_M54_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M54_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_209), .A2(
        top_AND_M54_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M54_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M54_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_306), .A2(top_AND_M54_U1_t_reg[5]), .ZN(
        top_AND_M54_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M54_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_210), .A2(
        top_AND_M54_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M54_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M54_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_305), .A2(top_AND_M54_U1_t_reg[6]), .ZN(
        top_AND_M54_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M54_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_209), .A2(
        top_AND_M54_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M54_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M54_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_305), .A2(top_AND_M54_U1_t_reg[7]), .ZN(
        top_AND_M54_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M54_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M54_U1_OperationInst_q[5]), .A2(
        top_AND_M54_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_338) );
  OR2_X1 top_AND_M54_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M54_U1_OperationInst_q[4]), .A2(
        top_AND_M54_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M54_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M54_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M54_U1_OperationInst_q[7]), .A2(
        top_AND_M54_U1_OperationInst_q[6]), .ZN(
        top_AND_M54_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M55_U1_nonlinearInst_U26 ( .A(top_AND_M55_U1_t[3]), .ZN(
        top_AND_M55_U1_t[7]) );
  OR2_X1 top_AND_M55_U1_nonlinearInst_U25 ( .A1(
        top_AND_M55_U1_nonlinearInst_n64), .A2(
        top_AND_M55_U1_nonlinearInst_n63), .ZN(top_AND_M55_U1_t[3]) );
  INV_X1 top_AND_M55_U1_nonlinearInst_U24 ( .A(
        top_AND_M55_U1_nonlinearInst_n62), .ZN(
        top_AND_M55_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M55_U1_nonlinearInst_U23 ( .A1(
        top_AND_M55_U1_nonlinearInst_n61), .A2(Fresh[25]), .ZN(
        top_AND_M55_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M55_U1_nonlinearInst_U22 ( .A1(Fresh[25]), .A2(
        top_AND_M55_U1_nonlinearInst_n61), .ZN(
        top_AND_M55_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M55_U1_nonlinearInst_U21 ( .A1(top_M44), .A2(top_T13), .ZN(
        top_AND_M55_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M55_U1_nonlinearInst_U20 ( .A(top_AND_M55_U1_t[2]), .ZN(
        top_AND_M55_U1_t[6]) );
  OR2_X1 top_AND_M55_U1_nonlinearInst_U19 ( .A1(
        top_AND_M55_U1_nonlinearInst_n60), .A2(
        top_AND_M55_U1_nonlinearInst_n59), .ZN(top_AND_M55_U1_t[2]) );
  INV_X1 top_AND_M55_U1_nonlinearInst_U18 ( .A(
        top_AND_M55_U1_nonlinearInst_n58), .ZN(
        top_AND_M55_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M55_U1_nonlinearInst_U17 ( .A1(
        top_AND_M55_U1_nonlinearInst_n57), .A2(Fresh[25]), .ZN(
        top_AND_M55_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M55_U1_nonlinearInst_U16 ( .A1(Fresh[25]), .A2(
        top_AND_M55_U1_nonlinearInst_n57), .ZN(
        top_AND_M55_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M55_U1_nonlinearInst_U15 ( .A1(
        top_AND_M55_U1_nonlinearInst_n56), .A2(top_M44), .ZN(
        top_AND_M55_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M55_U1_nonlinearInst_U14 ( .A(top_AND_M55_U1_t[1]), .ZN(
        top_AND_M55_U1_t[5]) );
  OR2_X1 top_AND_M55_U1_nonlinearInst_U13 ( .A1(
        top_AND_M55_U1_nonlinearInst_n55), .A2(
        top_AND_M55_U1_nonlinearInst_n54), .ZN(top_AND_M55_U1_t[1]) );
  AND2_X1 top_AND_M55_U1_nonlinearInst_U12 ( .A1(
        top_AND_M55_U1_nonlinearInst_n53), .A2(
        top_AND_M55_U1_nonlinearInst_n52), .ZN(
        top_AND_M55_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M55_U1_nonlinearInst_U11 ( .A(
        top_AND_M55_U1_nonlinearInst_n51), .ZN(
        top_AND_M55_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M55_U1_nonlinearInst_U10 ( .A1(
        top_AND_M55_U1_nonlinearInst_n52), .A2(
        top_AND_M55_U1_nonlinearInst_n53), .ZN(
        top_AND_M55_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M55_U1_nonlinearInst_U9 ( .A1(top_M44), .A2(
        top_AND_M55_U1_nonlinearInst_n56), .ZN(
        top_AND_M55_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M55_U1_nonlinearInst_U8 ( .A(top_T13), .ZN(
        top_AND_M55_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M55_U1_nonlinearInst_U7 ( .A(top_AND_M55_U1_t[0]), .ZN(
        top_AND_M55_U1_t[4]) );
  OR2_X1 top_AND_M55_U1_nonlinearInst_U6 ( .A1(
        top_AND_M55_U1_nonlinearInst_n50), .A2(
        top_AND_M55_U1_nonlinearInst_n49), .ZN(top_AND_M55_U1_t[0]) );
  AND2_X1 top_AND_M55_U1_nonlinearInst_U5 ( .A1(
        top_AND_M55_U1_nonlinearInst_n48), .A2(
        top_AND_M55_U1_nonlinearInst_n52), .ZN(
        top_AND_M55_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M55_U1_nonlinearInst_U4 ( .A(top_AND_M55_U1_nonlinearInst_n47), .ZN(top_AND_M55_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M55_U1_nonlinearInst_U3 ( .A1(
        top_AND_M55_U1_nonlinearInst_n52), .A2(
        top_AND_M55_U1_nonlinearInst_n48), .ZN(
        top_AND_M55_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M55_U1_nonlinearInst_U2 ( .A1(top_M44), .A2(top_T13), .ZN(
        top_AND_M55_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M55_U1_nonlinearInst_U1 ( .A(Fresh[25]), .ZN(
        top_AND_M55_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M55_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M55_U1_t[0]), .A2(
        top_AND_M55_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M55_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M55_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M55_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M55_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M55_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M55_U1_t_reg[0]) );
  AND2_X1 top_AND_M55_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M55_U1_t[1]), .A2(
        top_AND_M55_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M55_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M55_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M55_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M55_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M55_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M55_U1_t_reg[1]) );
  AND2_X1 top_AND_M55_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M55_U1_t[2]), .A2(
        top_AND_M55_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M55_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M55_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M55_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M55_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M55_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M55_U1_t_reg[2]) );
  AND2_X1 top_AND_M55_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M55_U1_t[3]), .A2(
        top_AND_M55_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M55_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M55_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M55_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M55_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M55_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M55_U1_t_reg[3]) );
  AND2_X1 top_AND_M55_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M55_U1_t[4]), .A2(
        top_AND_M55_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M55_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M55_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M55_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M55_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M55_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M55_U1_t_reg[4]) );
  AND2_X1 top_AND_M55_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M55_U1_t[5]), .A2(
        top_AND_M55_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M55_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M55_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M55_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M55_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M55_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M55_U1_t_reg[5]) );
  AND2_X1 top_AND_M55_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M55_U1_t[6]), .A2(
        top_AND_M55_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M55_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M55_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M55_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M55_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M55_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M55_U1_t_reg[6]) );
  AND2_X1 top_AND_M55_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M55_U1_t[7]), .A2(
        top_AND_M55_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M55_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M55_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M55_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M55_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M55_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M55_U1_t_reg[7]) );
  AND2_X1 top_AND_M55_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_196), .A2(
        top_AND_M55_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M55_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M55_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_312), .A2(top_AND_M55_U1_t_reg[0]), .ZN(
        top_AND_M55_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M55_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_195), .A2(
        top_AND_M55_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M55_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M55_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_312), .A2(top_AND_M55_U1_t_reg[1]), .ZN(
        top_AND_M55_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M55_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_196), .A2(
        top_AND_M55_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M55_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M55_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_311), .A2(top_AND_M55_U1_t_reg[2]), .ZN(
        top_AND_M55_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M55_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_195), .A2(
        top_AND_M55_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M55_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M55_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_311), .A2(top_AND_M55_U1_t_reg[3]), .ZN(
        top_AND_M55_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M55_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M55_U1_OperationInst_q[1]), .A2(
        top_AND_M55_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_339) );
  OR2_X1 top_AND_M55_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M55_U1_OperationInst_q[0]), .A2(
        top_AND_M55_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M55_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M55_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M55_U1_OperationInst_q[3]), .A2(
        top_AND_M55_U1_OperationInst_q[2]), .ZN(
        top_AND_M55_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M55_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_196), .A2(
        top_AND_M55_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M55_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M55_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_312), .A2(top_AND_M55_U1_t_reg[4]), .ZN(
        top_AND_M55_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M55_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_195), .A2(
        top_AND_M55_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M55_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M55_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_312), .A2(top_AND_M55_U1_t_reg[5]), .ZN(
        top_AND_M55_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M55_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_196), .A2(
        top_AND_M55_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M55_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M55_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_311), .A2(top_AND_M55_U1_t_reg[6]), .ZN(
        top_AND_M55_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M55_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_195), .A2(
        top_AND_M55_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M55_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M55_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_311), .A2(top_AND_M55_U1_t_reg[7]), .ZN(
        top_AND_M55_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M55_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M55_U1_OperationInst_q[5]), .A2(
        top_AND_M55_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_340) );
  OR2_X1 top_AND_M55_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M55_U1_OperationInst_q[4]), .A2(
        top_AND_M55_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M55_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M55_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M55_U1_OperationInst_q[7]), .A2(
        top_AND_M55_U1_OperationInst_q[6]), .ZN(
        top_AND_M55_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M56_U1_nonlinearInst_U26 ( .A(top_AND_M56_U1_t[0]), .ZN(
        top_AND_M56_U1_t[4]) );
  OR2_X1 top_AND_M56_U1_nonlinearInst_U25 ( .A1(
        top_AND_M56_U1_nonlinearInst_n64), .A2(
        top_AND_M56_U1_nonlinearInst_n63), .ZN(top_AND_M56_U1_t[0]) );
  AND2_X1 top_AND_M56_U1_nonlinearInst_U24 ( .A1(
        top_AND_M56_U1_nonlinearInst_n62), .A2(
        top_AND_M56_U1_nonlinearInst_n61), .ZN(
        top_AND_M56_U1_nonlinearInst_n63) );
  INV_X1 top_AND_M56_U1_nonlinearInst_U23 ( .A(
        top_AND_M56_U1_nonlinearInst_n60), .ZN(
        top_AND_M56_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M56_U1_nonlinearInst_U22 ( .A1(
        top_AND_M56_U1_nonlinearInst_n61), .A2(
        top_AND_M56_U1_nonlinearInst_n62), .ZN(
        top_AND_M56_U1_nonlinearInst_n60) );
  AND2_X1 top_AND_M56_U1_nonlinearInst_U21 ( .A1(top_M40), .A2(top_T23), .ZN(
        top_AND_M56_U1_nonlinearInst_n62) );
  INV_X1 top_AND_M56_U1_nonlinearInst_U20 ( .A(top_AND_M56_U1_t[3]), .ZN(
        top_AND_M56_U1_t[7]) );
  OR2_X1 top_AND_M56_U1_nonlinearInst_U19 ( .A1(
        top_AND_M56_U1_nonlinearInst_n59), .A2(
        top_AND_M56_U1_nonlinearInst_n58), .ZN(top_AND_M56_U1_t[3]) );
  INV_X1 top_AND_M56_U1_nonlinearInst_U18 ( .A(
        top_AND_M56_U1_nonlinearInst_n57), .ZN(
        top_AND_M56_U1_nonlinearInst_n58) );
  OR2_X1 top_AND_M56_U1_nonlinearInst_U17 ( .A1(
        top_AND_M56_U1_nonlinearInst_n56), .A2(Fresh[26]), .ZN(
        top_AND_M56_U1_nonlinearInst_n57) );
  AND2_X1 top_AND_M56_U1_nonlinearInst_U16 ( .A1(Fresh[26]), .A2(
        top_AND_M56_U1_nonlinearInst_n56), .ZN(
        top_AND_M56_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M56_U1_nonlinearInst_U15 ( .A1(top_M40), .A2(top_T23), .ZN(
        top_AND_M56_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M56_U1_nonlinearInst_U14 ( .A(top_AND_M56_U1_t[2]), .ZN(
        top_AND_M56_U1_t[6]) );
  OR2_X1 top_AND_M56_U1_nonlinearInst_U13 ( .A1(
        top_AND_M56_U1_nonlinearInst_n55), .A2(
        top_AND_M56_U1_nonlinearInst_n54), .ZN(top_AND_M56_U1_t[2]) );
  INV_X1 top_AND_M56_U1_nonlinearInst_U12 ( .A(
        top_AND_M56_U1_nonlinearInst_n53), .ZN(
        top_AND_M56_U1_nonlinearInst_n54) );
  OR2_X1 top_AND_M56_U1_nonlinearInst_U11 ( .A1(
        top_AND_M56_U1_nonlinearInst_n52), .A2(Fresh[26]), .ZN(
        top_AND_M56_U1_nonlinearInst_n53) );
  AND2_X1 top_AND_M56_U1_nonlinearInst_U10 ( .A1(Fresh[26]), .A2(
        top_AND_M56_U1_nonlinearInst_n52), .ZN(
        top_AND_M56_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M56_U1_nonlinearInst_U9 ( .A1(
        top_AND_M56_U1_nonlinearInst_n51), .A2(top_M40), .ZN(
        top_AND_M56_U1_nonlinearInst_n52) );
  INV_X1 top_AND_M56_U1_nonlinearInst_U8 ( .A(top_AND_M56_U1_t[1]), .ZN(
        top_AND_M56_U1_t[5]) );
  OR2_X1 top_AND_M56_U1_nonlinearInst_U7 ( .A1(
        top_AND_M56_U1_nonlinearInst_n50), .A2(
        top_AND_M56_U1_nonlinearInst_n49), .ZN(top_AND_M56_U1_t[1]) );
  AND2_X1 top_AND_M56_U1_nonlinearInst_U6 ( .A1(
        top_AND_M56_U1_nonlinearInst_n48), .A2(
        top_AND_M56_U1_nonlinearInst_n61), .ZN(
        top_AND_M56_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M56_U1_nonlinearInst_U5 ( .A(top_AND_M56_U1_nonlinearInst_n47), .ZN(top_AND_M56_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M56_U1_nonlinearInst_U4 ( .A1(
        top_AND_M56_U1_nonlinearInst_n61), .A2(
        top_AND_M56_U1_nonlinearInst_n48), .ZN(
        top_AND_M56_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M56_U1_nonlinearInst_U3 ( .A1(top_M40), .A2(
        top_AND_M56_U1_nonlinearInst_n51), .ZN(
        top_AND_M56_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M56_U1_nonlinearInst_U2 ( .A(top_T23), .ZN(
        top_AND_M56_U1_nonlinearInst_n51) );
  INV_X1 top_AND_M56_U1_nonlinearInst_U1 ( .A(Fresh[26]), .ZN(
        top_AND_M56_U1_nonlinearInst_n61) );
  AND2_X1 top_AND_M56_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M56_U1_t[0]), .A2(
        top_AND_M56_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M56_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M56_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M56_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M56_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M56_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M56_U1_t_reg[0]) );
  AND2_X1 top_AND_M56_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M56_U1_t[1]), .A2(
        top_AND_M56_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M56_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M56_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M56_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M56_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M56_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M56_U1_t_reg[1]) );
  AND2_X1 top_AND_M56_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M56_U1_t[2]), .A2(
        top_AND_M56_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M56_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M56_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M56_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M56_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M56_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M56_U1_t_reg[2]) );
  AND2_X1 top_AND_M56_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M56_U1_t[3]), .A2(
        top_AND_M56_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M56_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M56_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M56_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M56_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M56_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M56_U1_t_reg[3]) );
  AND2_X1 top_AND_M56_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M56_U1_t[4]), .A2(
        top_AND_M56_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M56_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M56_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M56_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M56_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M56_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M56_U1_t_reg[4]) );
  AND2_X1 top_AND_M56_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M56_U1_t[5]), .A2(
        top_AND_M56_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M56_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M56_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M56_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M56_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M56_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M56_U1_t_reg[5]) );
  AND2_X1 top_AND_M56_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M56_U1_t[6]), .A2(
        top_AND_M56_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M56_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M56_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M56_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M56_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M56_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M56_U1_t_reg[6]) );
  AND2_X1 top_AND_M56_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M56_U1_t[7]), .A2(
        top_AND_M56_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M56_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M56_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M56_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M56_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M56_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M56_U1_t_reg[7]) );
  AND2_X1 top_AND_M56_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_218), .A2(
        top_AND_M56_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M56_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M56_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_304), .A2(top_AND_M56_U1_t_reg[0]), .ZN(
        top_AND_M56_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M56_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_217), .A2(
        top_AND_M56_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M56_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M56_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_304), .A2(top_AND_M56_U1_t_reg[1]), .ZN(
        top_AND_M56_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M56_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_218), .A2(
        top_AND_M56_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M56_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M56_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_303), .A2(top_AND_M56_U1_t_reg[2]), .ZN(
        top_AND_M56_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M56_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_217), .A2(
        top_AND_M56_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M56_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M56_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_303), .A2(top_AND_M56_U1_t_reg[3]), .ZN(
        top_AND_M56_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M56_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M56_U1_OperationInst_q[1]), .A2(
        top_AND_M56_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_321) );
  OR2_X1 top_AND_M56_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M56_U1_OperationInst_q[0]), .A2(
        top_AND_M56_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M56_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M56_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M56_U1_OperationInst_q[3]), .A2(
        top_AND_M56_U1_OperationInst_q[2]), .ZN(
        top_AND_M56_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M56_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_218), .A2(
        top_AND_M56_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M56_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M56_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_304), .A2(top_AND_M56_U1_t_reg[4]), .ZN(
        top_AND_M56_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M56_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_217), .A2(
        top_AND_M56_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M56_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M56_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_304), .A2(top_AND_M56_U1_t_reg[5]), .ZN(
        top_AND_M56_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M56_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_218), .A2(
        top_AND_M56_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M56_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M56_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_303), .A2(top_AND_M56_U1_t_reg[6]), .ZN(
        top_AND_M56_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M56_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_217), .A2(
        top_AND_M56_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M56_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M56_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_303), .A2(top_AND_M56_U1_t_reg[7]), .ZN(
        top_AND_M56_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M56_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M56_U1_OperationInst_q[5]), .A2(
        top_AND_M56_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_322) );
  OR2_X1 top_AND_M56_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M56_U1_OperationInst_q[4]), .A2(
        top_AND_M56_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M56_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M56_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M56_U1_OperationInst_q[7]), .A2(
        top_AND_M56_U1_OperationInst_q[6]), .ZN(
        top_AND_M56_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M57_U1_nonlinearInst_U26 ( .A(top_AND_M57_U1_t[3]), .ZN(
        top_AND_M57_U1_t[7]) );
  OR2_X1 top_AND_M57_U1_nonlinearInst_U25 ( .A1(
        top_AND_M57_U1_nonlinearInst_n64), .A2(
        top_AND_M57_U1_nonlinearInst_n63), .ZN(top_AND_M57_U1_t[3]) );
  INV_X1 top_AND_M57_U1_nonlinearInst_U24 ( .A(
        top_AND_M57_U1_nonlinearInst_n62), .ZN(
        top_AND_M57_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M57_U1_nonlinearInst_U23 ( .A1(
        top_AND_M57_U1_nonlinearInst_n61), .A2(Fresh[27]), .ZN(
        top_AND_M57_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M57_U1_nonlinearInst_U22 ( .A1(Fresh[27]), .A2(
        top_AND_M57_U1_nonlinearInst_n61), .ZN(
        top_AND_M57_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M57_U1_nonlinearInst_U21 ( .A1(top_M39), .A2(top_T19), .ZN(
        top_AND_M57_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M57_U1_nonlinearInst_U20 ( .A(top_AND_M57_U1_t[2]), .ZN(
        top_AND_M57_U1_t[6]) );
  OR2_X1 top_AND_M57_U1_nonlinearInst_U19 ( .A1(
        top_AND_M57_U1_nonlinearInst_n60), .A2(
        top_AND_M57_U1_nonlinearInst_n59), .ZN(top_AND_M57_U1_t[2]) );
  INV_X1 top_AND_M57_U1_nonlinearInst_U18 ( .A(
        top_AND_M57_U1_nonlinearInst_n58), .ZN(
        top_AND_M57_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M57_U1_nonlinearInst_U17 ( .A1(
        top_AND_M57_U1_nonlinearInst_n57), .A2(Fresh[27]), .ZN(
        top_AND_M57_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M57_U1_nonlinearInst_U16 ( .A1(Fresh[27]), .A2(
        top_AND_M57_U1_nonlinearInst_n57), .ZN(
        top_AND_M57_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M57_U1_nonlinearInst_U15 ( .A1(
        top_AND_M57_U1_nonlinearInst_n56), .A2(top_M39), .ZN(
        top_AND_M57_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M57_U1_nonlinearInst_U14 ( .A(top_AND_M57_U1_t[1]), .ZN(
        top_AND_M57_U1_t[5]) );
  OR2_X1 top_AND_M57_U1_nonlinearInst_U13 ( .A1(
        top_AND_M57_U1_nonlinearInst_n55), .A2(
        top_AND_M57_U1_nonlinearInst_n54), .ZN(top_AND_M57_U1_t[1]) );
  AND2_X1 top_AND_M57_U1_nonlinearInst_U12 ( .A1(
        top_AND_M57_U1_nonlinearInst_n53), .A2(
        top_AND_M57_U1_nonlinearInst_n52), .ZN(
        top_AND_M57_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M57_U1_nonlinearInst_U11 ( .A(
        top_AND_M57_U1_nonlinearInst_n51), .ZN(
        top_AND_M57_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M57_U1_nonlinearInst_U10 ( .A1(
        top_AND_M57_U1_nonlinearInst_n52), .A2(
        top_AND_M57_U1_nonlinearInst_n53), .ZN(
        top_AND_M57_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M57_U1_nonlinearInst_U9 ( .A1(top_M39), .A2(
        top_AND_M57_U1_nonlinearInst_n56), .ZN(
        top_AND_M57_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M57_U1_nonlinearInst_U8 ( .A(top_T19), .ZN(
        top_AND_M57_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M57_U1_nonlinearInst_U7 ( .A(top_AND_M57_U1_t[0]), .ZN(
        top_AND_M57_U1_t[4]) );
  OR2_X1 top_AND_M57_U1_nonlinearInst_U6 ( .A1(
        top_AND_M57_U1_nonlinearInst_n50), .A2(
        top_AND_M57_U1_nonlinearInst_n49), .ZN(top_AND_M57_U1_t[0]) );
  AND2_X1 top_AND_M57_U1_nonlinearInst_U5 ( .A1(
        top_AND_M57_U1_nonlinearInst_n48), .A2(
        top_AND_M57_U1_nonlinearInst_n52), .ZN(
        top_AND_M57_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M57_U1_nonlinearInst_U4 ( .A(top_AND_M57_U1_nonlinearInst_n47), .ZN(top_AND_M57_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M57_U1_nonlinearInst_U3 ( .A1(
        top_AND_M57_U1_nonlinearInst_n52), .A2(
        top_AND_M57_U1_nonlinearInst_n48), .ZN(
        top_AND_M57_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M57_U1_nonlinearInst_U2 ( .A1(top_M39), .A2(top_T19), .ZN(
        top_AND_M57_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M57_U1_nonlinearInst_U1 ( .A(Fresh[27]), .ZN(
        top_AND_M57_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M57_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M57_U1_t[0]), .A2(
        top_AND_M57_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M57_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M57_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M57_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M57_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M57_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M57_U1_t_reg[0]) );
  AND2_X1 top_AND_M57_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M57_U1_t[1]), .A2(
        top_AND_M57_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M57_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M57_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M57_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M57_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M57_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M57_U1_t_reg[1]) );
  AND2_X1 top_AND_M57_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M57_U1_t[2]), .A2(
        top_AND_M57_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M57_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M57_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M57_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M57_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M57_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M57_U1_t_reg[2]) );
  AND2_X1 top_AND_M57_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M57_U1_t[3]), .A2(
        top_AND_M57_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M57_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M57_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M57_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M57_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M57_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M57_U1_t_reg[3]) );
  AND2_X1 top_AND_M57_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M57_U1_t[4]), .A2(
        top_AND_M57_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M57_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M57_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M57_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M57_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M57_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M57_U1_t_reg[4]) );
  AND2_X1 top_AND_M57_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M57_U1_t[5]), .A2(
        top_AND_M57_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M57_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M57_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M57_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M57_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M57_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M57_U1_t_reg[5]) );
  AND2_X1 top_AND_M57_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M57_U1_t[6]), .A2(
        top_AND_M57_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M57_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M57_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M57_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M57_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M57_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M57_U1_t_reg[6]) );
  AND2_X1 top_AND_M57_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M57_U1_t[7]), .A2(
        top_AND_M57_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M57_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M57_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M57_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M57_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M57_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M57_U1_t_reg[7]) );
  AND2_X1 top_AND_M57_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_202), .A2(
        top_AND_M57_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M57_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M57_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_302), .A2(top_AND_M57_U1_t_reg[0]), .ZN(
        top_AND_M57_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M57_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_201), .A2(
        top_AND_M57_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M57_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M57_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_302), .A2(top_AND_M57_U1_t_reg[1]), .ZN(
        top_AND_M57_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M57_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_202), .A2(
        top_AND_M57_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M57_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M57_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_301), .A2(top_AND_M57_U1_t_reg[2]), .ZN(
        top_AND_M57_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M57_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_201), .A2(
        top_AND_M57_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M57_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M57_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_301), .A2(top_AND_M57_U1_t_reg[3]), .ZN(
        top_AND_M57_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M57_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M57_U1_OperationInst_q[1]), .A2(
        top_AND_M57_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_323) );
  OR2_X1 top_AND_M57_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M57_U1_OperationInst_q[0]), .A2(
        top_AND_M57_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M57_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M57_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M57_U1_OperationInst_q[3]), .A2(
        top_AND_M57_U1_OperationInst_q[2]), .ZN(
        top_AND_M57_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M57_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_202), .A2(
        top_AND_M57_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M57_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M57_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_302), .A2(top_AND_M57_U1_t_reg[4]), .ZN(
        top_AND_M57_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M57_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_201), .A2(
        top_AND_M57_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M57_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M57_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_302), .A2(top_AND_M57_U1_t_reg[5]), .ZN(
        top_AND_M57_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M57_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_202), .A2(
        top_AND_M57_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M57_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M57_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_301), .A2(top_AND_M57_U1_t_reg[6]), .ZN(
        top_AND_M57_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M57_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_201), .A2(
        top_AND_M57_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M57_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M57_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_301), .A2(top_AND_M57_U1_t_reg[7]), .ZN(
        top_AND_M57_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M57_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M57_U1_OperationInst_q[5]), .A2(
        top_AND_M57_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_324) );
  OR2_X1 top_AND_M57_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M57_U1_OperationInst_q[4]), .A2(
        top_AND_M57_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M57_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M57_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M57_U1_OperationInst_q[7]), .A2(
        top_AND_M57_U1_OperationInst_q[6]), .ZN(
        top_AND_M57_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M58_U1_nonlinearInst_U26 ( .A(top_AND_M58_U1_t[3]), .ZN(
        top_AND_M58_U1_t[7]) );
  OR2_X1 top_AND_M58_U1_nonlinearInst_U25 ( .A1(
        top_AND_M58_U1_nonlinearInst_n64), .A2(
        top_AND_M58_U1_nonlinearInst_n63), .ZN(top_AND_M58_U1_t[3]) );
  INV_X1 top_AND_M58_U1_nonlinearInst_U24 ( .A(
        top_AND_M58_U1_nonlinearInst_n62), .ZN(
        top_AND_M58_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M58_U1_nonlinearInst_U23 ( .A1(
        top_AND_M58_U1_nonlinearInst_n61), .A2(Fresh[28]), .ZN(
        top_AND_M58_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M58_U1_nonlinearInst_U22 ( .A1(Fresh[28]), .A2(
        top_AND_M58_U1_nonlinearInst_n61), .ZN(
        top_AND_M58_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M58_U1_nonlinearInst_U21 ( .A1(top_M43), .A2(top_T3), .ZN(
        top_AND_M58_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M58_U1_nonlinearInst_U20 ( .A(top_AND_M58_U1_t[2]), .ZN(
        top_AND_M58_U1_t[6]) );
  OR2_X1 top_AND_M58_U1_nonlinearInst_U19 ( .A1(
        top_AND_M58_U1_nonlinearInst_n60), .A2(
        top_AND_M58_U1_nonlinearInst_n59), .ZN(top_AND_M58_U1_t[2]) );
  INV_X1 top_AND_M58_U1_nonlinearInst_U18 ( .A(
        top_AND_M58_U1_nonlinearInst_n58), .ZN(
        top_AND_M58_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M58_U1_nonlinearInst_U17 ( .A1(
        top_AND_M58_U1_nonlinearInst_n57), .A2(Fresh[28]), .ZN(
        top_AND_M58_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M58_U1_nonlinearInst_U16 ( .A1(Fresh[28]), .A2(
        top_AND_M58_U1_nonlinearInst_n57), .ZN(
        top_AND_M58_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M58_U1_nonlinearInst_U15 ( .A1(
        top_AND_M58_U1_nonlinearInst_n56), .A2(top_M43), .ZN(
        top_AND_M58_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M58_U1_nonlinearInst_U14 ( .A(top_AND_M58_U1_t[1]), .ZN(
        top_AND_M58_U1_t[5]) );
  OR2_X1 top_AND_M58_U1_nonlinearInst_U13 ( .A1(
        top_AND_M58_U1_nonlinearInst_n55), .A2(
        top_AND_M58_U1_nonlinearInst_n54), .ZN(top_AND_M58_U1_t[1]) );
  AND2_X1 top_AND_M58_U1_nonlinearInst_U12 ( .A1(
        top_AND_M58_U1_nonlinearInst_n53), .A2(
        top_AND_M58_U1_nonlinearInst_n52), .ZN(
        top_AND_M58_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M58_U1_nonlinearInst_U11 ( .A(
        top_AND_M58_U1_nonlinearInst_n51), .ZN(
        top_AND_M58_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M58_U1_nonlinearInst_U10 ( .A1(
        top_AND_M58_U1_nonlinearInst_n52), .A2(
        top_AND_M58_U1_nonlinearInst_n53), .ZN(
        top_AND_M58_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M58_U1_nonlinearInst_U9 ( .A1(top_M43), .A2(
        top_AND_M58_U1_nonlinearInst_n56), .ZN(
        top_AND_M58_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M58_U1_nonlinearInst_U8 ( .A(top_T3), .ZN(
        top_AND_M58_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M58_U1_nonlinearInst_U7 ( .A(top_AND_M58_U1_t[0]), .ZN(
        top_AND_M58_U1_t[4]) );
  OR2_X1 top_AND_M58_U1_nonlinearInst_U6 ( .A1(
        top_AND_M58_U1_nonlinearInst_n50), .A2(
        top_AND_M58_U1_nonlinearInst_n49), .ZN(top_AND_M58_U1_t[0]) );
  AND2_X1 top_AND_M58_U1_nonlinearInst_U5 ( .A1(
        top_AND_M58_U1_nonlinearInst_n48), .A2(
        top_AND_M58_U1_nonlinearInst_n52), .ZN(
        top_AND_M58_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M58_U1_nonlinearInst_U4 ( .A(top_AND_M58_U1_nonlinearInst_n47), .ZN(top_AND_M58_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M58_U1_nonlinearInst_U3 ( .A1(
        top_AND_M58_U1_nonlinearInst_n52), .A2(
        top_AND_M58_U1_nonlinearInst_n48), .ZN(
        top_AND_M58_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M58_U1_nonlinearInst_U2 ( .A1(top_M43), .A2(top_T3), .ZN(
        top_AND_M58_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M58_U1_nonlinearInst_U1 ( .A(Fresh[28]), .ZN(
        top_AND_M58_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M58_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M58_U1_t[0]), .A2(
        top_AND_M58_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M58_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M58_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M58_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M58_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M58_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M58_U1_t_reg[0]) );
  AND2_X1 top_AND_M58_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M58_U1_t[1]), .A2(
        top_AND_M58_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M58_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M58_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M58_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M58_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M58_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M58_U1_t_reg[1]) );
  AND2_X1 top_AND_M58_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M58_U1_t[2]), .A2(
        top_AND_M58_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M58_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M58_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M58_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M58_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M58_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M58_U1_t_reg[2]) );
  AND2_X1 top_AND_M58_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M58_U1_t[3]), .A2(
        top_AND_M58_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M58_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M58_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M58_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M58_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M58_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M58_U1_t_reg[3]) );
  AND2_X1 top_AND_M58_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M58_U1_t[4]), .A2(
        top_AND_M58_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M58_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M58_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M58_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M58_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M58_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M58_U1_t_reg[4]) );
  AND2_X1 top_AND_M58_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M58_U1_t[5]), .A2(
        top_AND_M58_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M58_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M58_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M58_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M58_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M58_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M58_U1_t_reg[5]) );
  AND2_X1 top_AND_M58_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M58_U1_t[6]), .A2(
        top_AND_M58_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M58_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M58_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M58_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M58_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M58_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M58_U1_t_reg[6]) );
  AND2_X1 top_AND_M58_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M58_U1_t[7]), .A2(
        top_AND_M58_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M58_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M58_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M58_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M58_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M58_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M58_U1_t_reg[7]) );
  AND2_X1 top_AND_M58_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_168), .A2(
        top_AND_M58_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M58_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M58_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_310), .A2(top_AND_M58_U1_t_reg[0]), .ZN(
        top_AND_M58_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M58_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_167), .A2(
        top_AND_M58_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M58_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M58_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_310), .A2(top_AND_M58_U1_t_reg[1]), .ZN(
        top_AND_M58_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M58_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_168), .A2(
        top_AND_M58_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M58_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M58_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_309), .A2(top_AND_M58_U1_t_reg[2]), .ZN(
        top_AND_M58_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M58_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_167), .A2(
        top_AND_M58_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M58_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M58_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_309), .A2(top_AND_M58_U1_t_reg[3]), .ZN(
        top_AND_M58_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M58_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M58_U1_OperationInst_q[1]), .A2(
        top_AND_M58_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_341) );
  OR2_X1 top_AND_M58_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M58_U1_OperationInst_q[0]), .A2(
        top_AND_M58_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M58_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M58_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M58_U1_OperationInst_q[3]), .A2(
        top_AND_M58_U1_OperationInst_q[2]), .ZN(
        top_AND_M58_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M58_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_168), .A2(
        top_AND_M58_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M58_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M58_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_310), .A2(top_AND_M58_U1_t_reg[4]), .ZN(
        top_AND_M58_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M58_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_167), .A2(
        top_AND_M58_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M58_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M58_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_310), .A2(top_AND_M58_U1_t_reg[5]), .ZN(
        top_AND_M58_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M58_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_168), .A2(
        top_AND_M58_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M58_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M58_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_309), .A2(top_AND_M58_U1_t_reg[6]), .ZN(
        top_AND_M58_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M58_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_167), .A2(
        top_AND_M58_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M58_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M58_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_309), .A2(top_AND_M58_U1_t_reg[7]), .ZN(
        top_AND_M58_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M58_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M58_U1_OperationInst_q[5]), .A2(
        top_AND_M58_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_342) );
  OR2_X1 top_AND_M58_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M58_U1_OperationInst_q[4]), .A2(
        top_AND_M58_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M58_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M58_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M58_U1_OperationInst_q[7]), .A2(
        top_AND_M58_U1_OperationInst_q[6]), .ZN(
        top_AND_M58_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M59_U1_nonlinearInst_U26 ( .A(top_AND_M59_U1_t[3]), .ZN(
        top_AND_M59_U1_t[7]) );
  OR2_X1 top_AND_M59_U1_nonlinearInst_U25 ( .A1(
        top_AND_M59_U1_nonlinearInst_n64), .A2(
        top_AND_M59_U1_nonlinearInst_n63), .ZN(top_AND_M59_U1_t[3]) );
  INV_X1 top_AND_M59_U1_nonlinearInst_U24 ( .A(
        top_AND_M59_U1_nonlinearInst_n62), .ZN(
        top_AND_M59_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M59_U1_nonlinearInst_U23 ( .A1(
        top_AND_M59_U1_nonlinearInst_n61), .A2(Fresh[29]), .ZN(
        top_AND_M59_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M59_U1_nonlinearInst_U22 ( .A1(Fresh[29]), .A2(
        top_AND_M59_U1_nonlinearInst_n61), .ZN(
        top_AND_M59_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M59_U1_nonlinearInst_U21 ( .A1(top_M38), .A2(top_T22), .ZN(
        top_AND_M59_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M59_U1_nonlinearInst_U20 ( .A(top_AND_M59_U1_t[2]), .ZN(
        top_AND_M59_U1_t[6]) );
  OR2_X1 top_AND_M59_U1_nonlinearInst_U19 ( .A1(
        top_AND_M59_U1_nonlinearInst_n60), .A2(
        top_AND_M59_U1_nonlinearInst_n59), .ZN(top_AND_M59_U1_t[2]) );
  INV_X1 top_AND_M59_U1_nonlinearInst_U18 ( .A(
        top_AND_M59_U1_nonlinearInst_n58), .ZN(
        top_AND_M59_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M59_U1_nonlinearInst_U17 ( .A1(
        top_AND_M59_U1_nonlinearInst_n57), .A2(Fresh[29]), .ZN(
        top_AND_M59_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M59_U1_nonlinearInst_U16 ( .A1(Fresh[29]), .A2(
        top_AND_M59_U1_nonlinearInst_n57), .ZN(
        top_AND_M59_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M59_U1_nonlinearInst_U15 ( .A1(
        top_AND_M59_U1_nonlinearInst_n56), .A2(top_M38), .ZN(
        top_AND_M59_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M59_U1_nonlinearInst_U14 ( .A(top_AND_M59_U1_t[1]), .ZN(
        top_AND_M59_U1_t[5]) );
  OR2_X1 top_AND_M59_U1_nonlinearInst_U13 ( .A1(
        top_AND_M59_U1_nonlinearInst_n55), .A2(
        top_AND_M59_U1_nonlinearInst_n54), .ZN(top_AND_M59_U1_t[1]) );
  AND2_X1 top_AND_M59_U1_nonlinearInst_U12 ( .A1(
        top_AND_M59_U1_nonlinearInst_n53), .A2(
        top_AND_M59_U1_nonlinearInst_n52), .ZN(
        top_AND_M59_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M59_U1_nonlinearInst_U11 ( .A(
        top_AND_M59_U1_nonlinearInst_n51), .ZN(
        top_AND_M59_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M59_U1_nonlinearInst_U10 ( .A1(
        top_AND_M59_U1_nonlinearInst_n52), .A2(
        top_AND_M59_U1_nonlinearInst_n53), .ZN(
        top_AND_M59_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M59_U1_nonlinearInst_U9 ( .A1(top_M38), .A2(
        top_AND_M59_U1_nonlinearInst_n56), .ZN(
        top_AND_M59_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M59_U1_nonlinearInst_U8 ( .A(top_T22), .ZN(
        top_AND_M59_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M59_U1_nonlinearInst_U7 ( .A(top_AND_M59_U1_t[0]), .ZN(
        top_AND_M59_U1_t[4]) );
  OR2_X1 top_AND_M59_U1_nonlinearInst_U6 ( .A1(
        top_AND_M59_U1_nonlinearInst_n50), .A2(
        top_AND_M59_U1_nonlinearInst_n49), .ZN(top_AND_M59_U1_t[0]) );
  AND2_X1 top_AND_M59_U1_nonlinearInst_U5 ( .A1(
        top_AND_M59_U1_nonlinearInst_n48), .A2(
        top_AND_M59_U1_nonlinearInst_n52), .ZN(
        top_AND_M59_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M59_U1_nonlinearInst_U4 ( .A(top_AND_M59_U1_nonlinearInst_n47), .ZN(top_AND_M59_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M59_U1_nonlinearInst_U3 ( .A1(
        top_AND_M59_U1_nonlinearInst_n52), .A2(
        top_AND_M59_U1_nonlinearInst_n48), .ZN(
        top_AND_M59_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M59_U1_nonlinearInst_U2 ( .A1(top_M38), .A2(top_T22), .ZN(
        top_AND_M59_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M59_U1_nonlinearInst_U1 ( .A(Fresh[29]), .ZN(
        top_AND_M59_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M59_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M59_U1_t[0]), .A2(
        top_AND_M59_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M59_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M59_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M59_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M59_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M59_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M59_U1_t_reg[0]) );
  AND2_X1 top_AND_M59_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M59_U1_t[1]), .A2(
        top_AND_M59_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M59_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M59_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M59_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M59_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M59_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M59_U1_t_reg[1]) );
  AND2_X1 top_AND_M59_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M59_U1_t[2]), .A2(
        top_AND_M59_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M59_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M59_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M59_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M59_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M59_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M59_U1_t_reg[2]) );
  AND2_X1 top_AND_M59_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M59_U1_t[3]), .A2(
        top_AND_M59_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M59_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M59_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M59_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M59_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M59_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M59_U1_t_reg[3]) );
  AND2_X1 top_AND_M59_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M59_U1_t[4]), .A2(
        top_AND_M59_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M59_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M59_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M59_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M59_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M59_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M59_U1_t_reg[4]) );
  AND2_X1 top_AND_M59_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M59_U1_t[5]), .A2(
        top_AND_M59_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M59_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M59_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M59_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M59_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M59_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M59_U1_t_reg[5]) );
  AND2_X1 top_AND_M59_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M59_U1_t[6]), .A2(
        top_AND_M59_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M59_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M59_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M59_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M59_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M59_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M59_U1_t_reg[6]) );
  AND2_X1 top_AND_M59_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M59_U1_t[7]), .A2(
        top_AND_M59_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M59_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M59_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M59_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M59_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M59_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M59_U1_t_reg[7]) );
  AND2_X1 top_AND_M59_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_204), .A2(
        top_AND_M59_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M59_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M59_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_300), .A2(top_AND_M59_U1_t_reg[0]), .ZN(
        top_AND_M59_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M59_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_203), .A2(
        top_AND_M59_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M59_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M59_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_300), .A2(top_AND_M59_U1_t_reg[1]), .ZN(
        top_AND_M59_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M59_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_204), .A2(
        top_AND_M59_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M59_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M59_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_299), .A2(top_AND_M59_U1_t_reg[2]), .ZN(
        top_AND_M59_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M59_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_203), .A2(
        top_AND_M59_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M59_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M59_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_299), .A2(top_AND_M59_U1_t_reg[3]), .ZN(
        top_AND_M59_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M59_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M59_U1_OperationInst_q[1]), .A2(
        top_AND_M59_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_325) );
  OR2_X1 top_AND_M59_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M59_U1_OperationInst_q[0]), .A2(
        top_AND_M59_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M59_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M59_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M59_U1_OperationInst_q[3]), .A2(
        top_AND_M59_U1_OperationInst_q[2]), .ZN(
        top_AND_M59_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M59_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_204), .A2(
        top_AND_M59_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M59_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M59_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_300), .A2(top_AND_M59_U1_t_reg[4]), .ZN(
        top_AND_M59_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M59_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_203), .A2(
        top_AND_M59_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M59_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M59_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_300), .A2(top_AND_M59_U1_t_reg[5]), .ZN(
        top_AND_M59_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M59_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_204), .A2(
        top_AND_M59_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M59_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M59_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_299), .A2(top_AND_M59_U1_t_reg[6]), .ZN(
        top_AND_M59_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M59_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_203), .A2(
        top_AND_M59_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M59_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M59_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_299), .A2(top_AND_M59_U1_t_reg[7]), .ZN(
        top_AND_M59_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M59_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M59_U1_OperationInst_q[5]), .A2(
        top_AND_M59_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_326) );
  OR2_X1 top_AND_M59_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M59_U1_OperationInst_q[4]), .A2(
        top_AND_M59_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M59_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M59_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M59_U1_OperationInst_q[7]), .A2(
        top_AND_M59_U1_OperationInst_q[6]), .ZN(
        top_AND_M59_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M60_U1_nonlinearInst_U26 ( .A(top_AND_M60_U1_t[3]), .ZN(
        top_AND_M60_U1_t[7]) );
  OR2_X1 top_AND_M60_U1_nonlinearInst_U25 ( .A1(
        top_AND_M60_U1_nonlinearInst_n64), .A2(
        top_AND_M60_U1_nonlinearInst_n63), .ZN(top_AND_M60_U1_t[3]) );
  INV_X1 top_AND_M60_U1_nonlinearInst_U24 ( .A(
        top_AND_M60_U1_nonlinearInst_n62), .ZN(
        top_AND_M60_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M60_U1_nonlinearInst_U23 ( .A1(
        top_AND_M60_U1_nonlinearInst_n61), .A2(Fresh[30]), .ZN(
        top_AND_M60_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M60_U1_nonlinearInst_U22 ( .A1(Fresh[30]), .A2(
        top_AND_M60_U1_nonlinearInst_n61), .ZN(
        top_AND_M60_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M60_U1_nonlinearInst_U21 ( .A1(top_M37), .A2(top_T20), .ZN(
        top_AND_M60_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M60_U1_nonlinearInst_U20 ( .A(top_AND_M60_U1_t[2]), .ZN(
        top_AND_M60_U1_t[6]) );
  OR2_X1 top_AND_M60_U1_nonlinearInst_U19 ( .A1(
        top_AND_M60_U1_nonlinearInst_n60), .A2(
        top_AND_M60_U1_nonlinearInst_n59), .ZN(top_AND_M60_U1_t[2]) );
  INV_X1 top_AND_M60_U1_nonlinearInst_U18 ( .A(
        top_AND_M60_U1_nonlinearInst_n58), .ZN(
        top_AND_M60_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M60_U1_nonlinearInst_U17 ( .A1(
        top_AND_M60_U1_nonlinearInst_n57), .A2(Fresh[30]), .ZN(
        top_AND_M60_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M60_U1_nonlinearInst_U16 ( .A1(Fresh[30]), .A2(
        top_AND_M60_U1_nonlinearInst_n57), .ZN(
        top_AND_M60_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M60_U1_nonlinearInst_U15 ( .A1(
        top_AND_M60_U1_nonlinearInst_n56), .A2(top_M37), .ZN(
        top_AND_M60_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M60_U1_nonlinearInst_U14 ( .A(top_AND_M60_U1_t[1]), .ZN(
        top_AND_M60_U1_t[5]) );
  OR2_X1 top_AND_M60_U1_nonlinearInst_U13 ( .A1(
        top_AND_M60_U1_nonlinearInst_n55), .A2(
        top_AND_M60_U1_nonlinearInst_n54), .ZN(top_AND_M60_U1_t[1]) );
  AND2_X1 top_AND_M60_U1_nonlinearInst_U12 ( .A1(
        top_AND_M60_U1_nonlinearInst_n53), .A2(
        top_AND_M60_U1_nonlinearInst_n52), .ZN(
        top_AND_M60_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M60_U1_nonlinearInst_U11 ( .A(
        top_AND_M60_U1_nonlinearInst_n51), .ZN(
        top_AND_M60_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M60_U1_nonlinearInst_U10 ( .A1(
        top_AND_M60_U1_nonlinearInst_n52), .A2(
        top_AND_M60_U1_nonlinearInst_n53), .ZN(
        top_AND_M60_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M60_U1_nonlinearInst_U9 ( .A1(top_M37), .A2(
        top_AND_M60_U1_nonlinearInst_n56), .ZN(
        top_AND_M60_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M60_U1_nonlinearInst_U8 ( .A(top_T20), .ZN(
        top_AND_M60_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M60_U1_nonlinearInst_U7 ( .A(top_AND_M60_U1_t[0]), .ZN(
        top_AND_M60_U1_t[4]) );
  OR2_X1 top_AND_M60_U1_nonlinearInst_U6 ( .A1(
        top_AND_M60_U1_nonlinearInst_n50), .A2(
        top_AND_M60_U1_nonlinearInst_n49), .ZN(top_AND_M60_U1_t[0]) );
  AND2_X1 top_AND_M60_U1_nonlinearInst_U5 ( .A1(
        top_AND_M60_U1_nonlinearInst_n48), .A2(
        top_AND_M60_U1_nonlinearInst_n52), .ZN(
        top_AND_M60_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M60_U1_nonlinearInst_U4 ( .A(top_AND_M60_U1_nonlinearInst_n47), .ZN(top_AND_M60_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M60_U1_nonlinearInst_U3 ( .A1(
        top_AND_M60_U1_nonlinearInst_n52), .A2(
        top_AND_M60_U1_nonlinearInst_n48), .ZN(
        top_AND_M60_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M60_U1_nonlinearInst_U2 ( .A1(top_M37), .A2(top_T20), .ZN(
        top_AND_M60_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M60_U1_nonlinearInst_U1 ( .A(Fresh[30]), .ZN(
        top_AND_M60_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M60_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M60_U1_t[0]), .A2(
        top_AND_M60_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M60_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M60_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M60_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M60_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M60_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M60_U1_t_reg[0]) );
  AND2_X1 top_AND_M60_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M60_U1_t[1]), .A2(
        top_AND_M60_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M60_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M60_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M60_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M60_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M60_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M60_U1_t_reg[1]) );
  AND2_X1 top_AND_M60_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M60_U1_t[2]), .A2(
        top_AND_M60_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M60_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M60_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M60_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M60_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M60_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M60_U1_t_reg[2]) );
  AND2_X1 top_AND_M60_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M60_U1_t[3]), .A2(
        top_AND_M60_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M60_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M60_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M60_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M60_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M60_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M60_U1_t_reg[3]) );
  AND2_X1 top_AND_M60_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M60_U1_t[4]), .A2(
        top_AND_M60_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M60_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M60_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M60_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M60_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M60_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M60_U1_t_reg[4]) );
  AND2_X1 top_AND_M60_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M60_U1_t[5]), .A2(
        top_AND_M60_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M60_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M60_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M60_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M60_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M60_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M60_U1_t_reg[5]) );
  AND2_X1 top_AND_M60_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M60_U1_t[6]), .A2(
        top_AND_M60_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M60_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M60_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M60_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M60_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M60_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M60_U1_t_reg[6]) );
  AND2_X1 top_AND_M60_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M60_U1_t[7]), .A2(
        top_AND_M60_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M60_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M60_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M60_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M60_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M60_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M60_U1_t_reg[7]) );
  AND2_X1 top_AND_M60_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_216), .A2(
        top_AND_M60_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M60_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M60_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_298), .A2(top_AND_M60_U1_t_reg[0]), .ZN(
        top_AND_M60_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M60_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_215), .A2(
        top_AND_M60_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M60_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M60_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_298), .A2(top_AND_M60_U1_t_reg[1]), .ZN(
        top_AND_M60_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M60_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_216), .A2(
        top_AND_M60_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M60_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M60_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_297), .A2(top_AND_M60_U1_t_reg[2]), .ZN(
        top_AND_M60_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M60_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_215), .A2(
        top_AND_M60_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M60_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M60_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_297), .A2(top_AND_M60_U1_t_reg[3]), .ZN(
        top_AND_M60_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M60_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M60_U1_OperationInst_q[1]), .A2(
        top_AND_M60_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_327) );
  OR2_X1 top_AND_M60_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M60_U1_OperationInst_q[0]), .A2(
        top_AND_M60_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M60_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M60_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M60_U1_OperationInst_q[3]), .A2(
        top_AND_M60_U1_OperationInst_q[2]), .ZN(
        top_AND_M60_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M60_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_216), .A2(
        top_AND_M60_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M60_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M60_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_298), .A2(top_AND_M60_U1_t_reg[4]), .ZN(
        top_AND_M60_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M60_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_215), .A2(
        top_AND_M60_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M60_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M60_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_298), .A2(top_AND_M60_U1_t_reg[5]), .ZN(
        top_AND_M60_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M60_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_216), .A2(
        top_AND_M60_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M60_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M60_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_297), .A2(top_AND_M60_U1_t_reg[6]), .ZN(
        top_AND_M60_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M60_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_215), .A2(
        top_AND_M60_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M60_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M60_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_297), .A2(top_AND_M60_U1_t_reg[7]), .ZN(
        top_AND_M60_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M60_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M60_U1_OperationInst_q[5]), .A2(
        top_AND_M60_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_328) );
  OR2_X1 top_AND_M60_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M60_U1_OperationInst_q[4]), .A2(
        top_AND_M60_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M60_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M60_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M60_U1_OperationInst_q[7]), .A2(
        top_AND_M60_U1_OperationInst_q[6]), .ZN(
        top_AND_M60_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M61_U1_nonlinearInst_U26 ( .A(top_AND_M61_U1_t[3]), .ZN(
        top_AND_M61_U1_t[7]) );
  OR2_X1 top_AND_M61_U1_nonlinearInst_U25 ( .A1(
        top_AND_M61_U1_nonlinearInst_n64), .A2(
        top_AND_M61_U1_nonlinearInst_n63), .ZN(top_AND_M61_U1_t[3]) );
  INV_X1 top_AND_M61_U1_nonlinearInst_U24 ( .A(
        top_AND_M61_U1_nonlinearInst_n62), .ZN(
        top_AND_M61_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M61_U1_nonlinearInst_U23 ( .A1(
        top_AND_M61_U1_nonlinearInst_n61), .A2(Fresh[31]), .ZN(
        top_AND_M61_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M61_U1_nonlinearInst_U22 ( .A1(Fresh[31]), .A2(
        top_AND_M61_U1_nonlinearInst_n61), .ZN(
        top_AND_M61_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M61_U1_nonlinearInst_U21 ( .A1(top_M42), .A2(top_T1), .ZN(
        top_AND_M61_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M61_U1_nonlinearInst_U20 ( .A(top_AND_M61_U1_t[2]), .ZN(
        top_AND_M61_U1_t[6]) );
  OR2_X1 top_AND_M61_U1_nonlinearInst_U19 ( .A1(
        top_AND_M61_U1_nonlinearInst_n60), .A2(
        top_AND_M61_U1_nonlinearInst_n59), .ZN(top_AND_M61_U1_t[2]) );
  INV_X1 top_AND_M61_U1_nonlinearInst_U18 ( .A(
        top_AND_M61_U1_nonlinearInst_n58), .ZN(
        top_AND_M61_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M61_U1_nonlinearInst_U17 ( .A1(
        top_AND_M61_U1_nonlinearInst_n57), .A2(Fresh[31]), .ZN(
        top_AND_M61_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M61_U1_nonlinearInst_U16 ( .A1(Fresh[31]), .A2(
        top_AND_M61_U1_nonlinearInst_n57), .ZN(
        top_AND_M61_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M61_U1_nonlinearInst_U15 ( .A1(
        top_AND_M61_U1_nonlinearInst_n56), .A2(top_M42), .ZN(
        top_AND_M61_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M61_U1_nonlinearInst_U14 ( .A(top_AND_M61_U1_t[1]), .ZN(
        top_AND_M61_U1_t[5]) );
  OR2_X1 top_AND_M61_U1_nonlinearInst_U13 ( .A1(
        top_AND_M61_U1_nonlinearInst_n55), .A2(
        top_AND_M61_U1_nonlinearInst_n54), .ZN(top_AND_M61_U1_t[1]) );
  AND2_X1 top_AND_M61_U1_nonlinearInst_U12 ( .A1(
        top_AND_M61_U1_nonlinearInst_n53), .A2(
        top_AND_M61_U1_nonlinearInst_n52), .ZN(
        top_AND_M61_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M61_U1_nonlinearInst_U11 ( .A(
        top_AND_M61_U1_nonlinearInst_n51), .ZN(
        top_AND_M61_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M61_U1_nonlinearInst_U10 ( .A1(
        top_AND_M61_U1_nonlinearInst_n52), .A2(
        top_AND_M61_U1_nonlinearInst_n53), .ZN(
        top_AND_M61_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M61_U1_nonlinearInst_U9 ( .A1(top_M42), .A2(
        top_AND_M61_U1_nonlinearInst_n56), .ZN(
        top_AND_M61_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M61_U1_nonlinearInst_U8 ( .A(top_T1), .ZN(
        top_AND_M61_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M61_U1_nonlinearInst_U7 ( .A(top_AND_M61_U1_t[0]), .ZN(
        top_AND_M61_U1_t[4]) );
  OR2_X1 top_AND_M61_U1_nonlinearInst_U6 ( .A1(
        top_AND_M61_U1_nonlinearInst_n50), .A2(
        top_AND_M61_U1_nonlinearInst_n49), .ZN(top_AND_M61_U1_t[0]) );
  AND2_X1 top_AND_M61_U1_nonlinearInst_U5 ( .A1(
        top_AND_M61_U1_nonlinearInst_n48), .A2(
        top_AND_M61_U1_nonlinearInst_n52), .ZN(
        top_AND_M61_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M61_U1_nonlinearInst_U4 ( .A(top_AND_M61_U1_nonlinearInst_n47), .ZN(top_AND_M61_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M61_U1_nonlinearInst_U3 ( .A1(
        top_AND_M61_U1_nonlinearInst_n52), .A2(
        top_AND_M61_U1_nonlinearInst_n48), .ZN(
        top_AND_M61_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M61_U1_nonlinearInst_U2 ( .A1(top_M42), .A2(top_T1), .ZN(
        top_AND_M61_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M61_U1_nonlinearInst_U1 ( .A(Fresh[31]), .ZN(
        top_AND_M61_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M61_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M61_U1_t[0]), .A2(
        top_AND_M61_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M61_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M61_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M61_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M61_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M61_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M61_U1_t_reg[0]) );
  AND2_X1 top_AND_M61_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M61_U1_t[1]), .A2(
        top_AND_M61_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M61_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M61_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M61_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M61_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M61_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M61_U1_t_reg[1]) );
  AND2_X1 top_AND_M61_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M61_U1_t[2]), .A2(
        top_AND_M61_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M61_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M61_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M61_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M61_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M61_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M61_U1_t_reg[2]) );
  AND2_X1 top_AND_M61_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M61_U1_t[3]), .A2(
        top_AND_M61_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M61_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M61_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M61_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M61_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M61_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M61_U1_t_reg[3]) );
  AND2_X1 top_AND_M61_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M61_U1_t[4]), .A2(
        top_AND_M61_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M61_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M61_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M61_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M61_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M61_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M61_U1_t_reg[4]) );
  AND2_X1 top_AND_M61_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M61_U1_t[5]), .A2(
        top_AND_M61_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M61_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M61_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M61_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M61_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M61_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M61_U1_t_reg[5]) );
  AND2_X1 top_AND_M61_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M61_U1_t[6]), .A2(
        top_AND_M61_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M61_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M61_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M61_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M61_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M61_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M61_U1_t_reg[6]) );
  AND2_X1 top_AND_M61_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M61_U1_t[7]), .A2(
        top_AND_M61_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M61_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M61_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M61_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M61_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M61_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M61_U1_t_reg[7]) );
  AND2_X1 top_AND_M61_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_160), .A2(
        top_AND_M61_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M61_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M61_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_308), .A2(top_AND_M61_U1_t_reg[0]), .ZN(
        top_AND_M61_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M61_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_159), .A2(
        top_AND_M61_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M61_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M61_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_308), .A2(top_AND_M61_U1_t_reg[1]), .ZN(
        top_AND_M61_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M61_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_160), .A2(
        top_AND_M61_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M61_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M61_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_307), .A2(top_AND_M61_U1_t_reg[2]), .ZN(
        top_AND_M61_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M61_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_159), .A2(
        top_AND_M61_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M61_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M61_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_307), .A2(top_AND_M61_U1_t_reg[3]), .ZN(
        top_AND_M61_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M61_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M61_U1_OperationInst_q[1]), .A2(
        top_AND_M61_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_343) );
  OR2_X1 top_AND_M61_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M61_U1_OperationInst_q[0]), .A2(
        top_AND_M61_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M61_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M61_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M61_U1_OperationInst_q[3]), .A2(
        top_AND_M61_U1_OperationInst_q[2]), .ZN(
        top_AND_M61_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M61_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_160), .A2(
        top_AND_M61_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M61_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M61_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_308), .A2(top_AND_M61_U1_t_reg[4]), .ZN(
        top_AND_M61_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M61_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_159), .A2(
        top_AND_M61_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M61_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M61_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_308), .A2(top_AND_M61_U1_t_reg[5]), .ZN(
        top_AND_M61_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M61_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_160), .A2(
        top_AND_M61_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M61_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M61_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_307), .A2(top_AND_M61_U1_t_reg[6]), .ZN(
        top_AND_M61_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M61_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_159), .A2(
        top_AND_M61_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M61_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M61_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_307), .A2(top_AND_M61_U1_t_reg[7]), .ZN(
        top_AND_M61_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M61_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M61_U1_OperationInst_q[5]), .A2(
        top_AND_M61_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_344) );
  OR2_X1 top_AND_M61_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M61_U1_OperationInst_q[4]), .A2(
        top_AND_M61_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M61_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M61_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M61_U1_OperationInst_q[7]), .A2(
        top_AND_M61_U1_OperationInst_q[6]), .ZN(
        top_AND_M61_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M62_U1_nonlinearInst_U26 ( .A(top_AND_M62_U1_t[3]), .ZN(
        top_AND_M62_U1_t[7]) );
  OR2_X1 top_AND_M62_U1_nonlinearInst_U25 ( .A1(
        top_AND_M62_U1_nonlinearInst_n64), .A2(
        top_AND_M62_U1_nonlinearInst_n63), .ZN(top_AND_M62_U1_t[3]) );
  INV_X1 top_AND_M62_U1_nonlinearInst_U24 ( .A(
        top_AND_M62_U1_nonlinearInst_n62), .ZN(
        top_AND_M62_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M62_U1_nonlinearInst_U23 ( .A1(
        top_AND_M62_U1_nonlinearInst_n61), .A2(Fresh[32]), .ZN(
        top_AND_M62_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M62_U1_nonlinearInst_U22 ( .A1(Fresh[32]), .A2(
        top_AND_M62_U1_nonlinearInst_n61), .ZN(
        top_AND_M62_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M62_U1_nonlinearInst_U21 ( .A1(top_M45), .A2(top_T4), .ZN(
        top_AND_M62_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M62_U1_nonlinearInst_U20 ( .A(top_AND_M62_U1_t[2]), .ZN(
        top_AND_M62_U1_t[6]) );
  OR2_X1 top_AND_M62_U1_nonlinearInst_U19 ( .A1(
        top_AND_M62_U1_nonlinearInst_n60), .A2(
        top_AND_M62_U1_nonlinearInst_n59), .ZN(top_AND_M62_U1_t[2]) );
  INV_X1 top_AND_M62_U1_nonlinearInst_U18 ( .A(
        top_AND_M62_U1_nonlinearInst_n58), .ZN(
        top_AND_M62_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M62_U1_nonlinearInst_U17 ( .A1(
        top_AND_M62_U1_nonlinearInst_n57), .A2(Fresh[32]), .ZN(
        top_AND_M62_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M62_U1_nonlinearInst_U16 ( .A1(Fresh[32]), .A2(
        top_AND_M62_U1_nonlinearInst_n57), .ZN(
        top_AND_M62_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M62_U1_nonlinearInst_U15 ( .A1(
        top_AND_M62_U1_nonlinearInst_n56), .A2(top_M45), .ZN(
        top_AND_M62_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M62_U1_nonlinearInst_U14 ( .A(top_AND_M62_U1_t[1]), .ZN(
        top_AND_M62_U1_t[5]) );
  OR2_X1 top_AND_M62_U1_nonlinearInst_U13 ( .A1(
        top_AND_M62_U1_nonlinearInst_n55), .A2(
        top_AND_M62_U1_nonlinearInst_n54), .ZN(top_AND_M62_U1_t[1]) );
  AND2_X1 top_AND_M62_U1_nonlinearInst_U12 ( .A1(
        top_AND_M62_U1_nonlinearInst_n53), .A2(
        top_AND_M62_U1_nonlinearInst_n52), .ZN(
        top_AND_M62_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M62_U1_nonlinearInst_U11 ( .A(
        top_AND_M62_U1_nonlinearInst_n51), .ZN(
        top_AND_M62_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M62_U1_nonlinearInst_U10 ( .A1(
        top_AND_M62_U1_nonlinearInst_n52), .A2(
        top_AND_M62_U1_nonlinearInst_n53), .ZN(
        top_AND_M62_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M62_U1_nonlinearInst_U9 ( .A1(top_M45), .A2(
        top_AND_M62_U1_nonlinearInst_n56), .ZN(
        top_AND_M62_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M62_U1_nonlinearInst_U8 ( .A(top_T4), .ZN(
        top_AND_M62_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M62_U1_nonlinearInst_U7 ( .A(top_AND_M62_U1_t[0]), .ZN(
        top_AND_M62_U1_t[4]) );
  OR2_X1 top_AND_M62_U1_nonlinearInst_U6 ( .A1(
        top_AND_M62_U1_nonlinearInst_n50), .A2(
        top_AND_M62_U1_nonlinearInst_n49), .ZN(top_AND_M62_U1_t[0]) );
  AND2_X1 top_AND_M62_U1_nonlinearInst_U5 ( .A1(
        top_AND_M62_U1_nonlinearInst_n48), .A2(
        top_AND_M62_U1_nonlinearInst_n52), .ZN(
        top_AND_M62_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M62_U1_nonlinearInst_U4 ( .A(top_AND_M62_U1_nonlinearInst_n47), .ZN(top_AND_M62_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M62_U1_nonlinearInst_U3 ( .A1(
        top_AND_M62_U1_nonlinearInst_n52), .A2(
        top_AND_M62_U1_nonlinearInst_n48), .ZN(
        top_AND_M62_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M62_U1_nonlinearInst_U2 ( .A1(top_M45), .A2(top_T4), .ZN(
        top_AND_M62_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M62_U1_nonlinearInst_U1 ( .A(Fresh[32]), .ZN(
        top_AND_M62_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M62_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M62_U1_t[0]), .A2(
        top_AND_M62_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M62_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M62_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M62_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M62_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M62_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M62_U1_t_reg[0]) );
  AND2_X1 top_AND_M62_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M62_U1_t[1]), .A2(
        top_AND_M62_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M62_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M62_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M62_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M62_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M62_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M62_U1_t_reg[1]) );
  AND2_X1 top_AND_M62_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M62_U1_t[2]), .A2(
        top_AND_M62_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M62_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M62_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M62_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M62_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M62_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M62_U1_t_reg[2]) );
  AND2_X1 top_AND_M62_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M62_U1_t[3]), .A2(
        top_AND_M62_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M62_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M62_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M62_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M62_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M62_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M62_U1_t_reg[3]) );
  AND2_X1 top_AND_M62_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M62_U1_t[4]), .A2(
        top_AND_M62_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M62_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M62_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M62_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M62_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M62_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M62_U1_t_reg[4]) );
  AND2_X1 top_AND_M62_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M62_U1_t[5]), .A2(
        top_AND_M62_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M62_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M62_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M62_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M62_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M62_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M62_U1_t_reg[5]) );
  AND2_X1 top_AND_M62_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M62_U1_t[6]), .A2(
        top_AND_M62_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M62_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M62_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M62_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M62_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M62_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M62_U1_t_reg[6]) );
  AND2_X1 top_AND_M62_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M62_U1_t[7]), .A2(
        top_AND_M62_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M62_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M62_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M62_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M62_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M62_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M62_U1_t_reg[7]) );
  AND2_X1 top_AND_M62_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_170), .A2(
        top_AND_M62_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M62_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M62_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_330), .A2(top_AND_M62_U1_t_reg[0]), .ZN(
        top_AND_M62_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M62_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_169), .A2(
        top_AND_M62_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M62_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M62_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_330), .A2(top_AND_M62_U1_t_reg[1]), .ZN(
        top_AND_M62_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M62_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_170), .A2(
        top_AND_M62_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M62_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M62_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_329), .A2(top_AND_M62_U1_t_reg[2]), .ZN(
        top_AND_M62_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M62_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_169), .A2(
        top_AND_M62_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M62_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M62_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_329), .A2(top_AND_M62_U1_t_reg[3]), .ZN(
        top_AND_M62_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M62_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M62_U1_OperationInst_q[1]), .A2(
        top_AND_M62_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_355) );
  OR2_X1 top_AND_M62_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M62_U1_OperationInst_q[0]), .A2(
        top_AND_M62_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M62_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M62_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M62_U1_OperationInst_q[3]), .A2(
        top_AND_M62_U1_OperationInst_q[2]), .ZN(
        top_AND_M62_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M62_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_170), .A2(
        top_AND_M62_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M62_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M62_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_330), .A2(top_AND_M62_U1_t_reg[4]), .ZN(
        top_AND_M62_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M62_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_169), .A2(
        top_AND_M62_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M62_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M62_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_330), .A2(top_AND_M62_U1_t_reg[5]), .ZN(
        top_AND_M62_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M62_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_170), .A2(
        top_AND_M62_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M62_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M62_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_329), .A2(top_AND_M62_U1_t_reg[6]), .ZN(
        top_AND_M62_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M62_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_169), .A2(
        top_AND_M62_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M62_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M62_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_329), .A2(top_AND_M62_U1_t_reg[7]), .ZN(
        top_AND_M62_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M62_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M62_U1_OperationInst_q[5]), .A2(
        top_AND_M62_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_356) );
  OR2_X1 top_AND_M62_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M62_U1_OperationInst_q[4]), .A2(
        top_AND_M62_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M62_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M62_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M62_U1_OperationInst_q[7]), .A2(
        top_AND_M62_U1_OperationInst_q[6]), .ZN(
        top_AND_M62_U1_OperationInst_orInst2_n5) );
  INV_X1 top_AND_M63_U1_nonlinearInst_U26 ( .A(top_AND_M63_U1_t[3]), .ZN(
        top_AND_M63_U1_t[7]) );
  OR2_X1 top_AND_M63_U1_nonlinearInst_U25 ( .A1(
        top_AND_M63_U1_nonlinearInst_n64), .A2(
        top_AND_M63_U1_nonlinearInst_n63), .ZN(top_AND_M63_U1_t[3]) );
  INV_X1 top_AND_M63_U1_nonlinearInst_U24 ( .A(
        top_AND_M63_U1_nonlinearInst_n62), .ZN(
        top_AND_M63_U1_nonlinearInst_n63) );
  OR2_X1 top_AND_M63_U1_nonlinearInst_U23 ( .A1(
        top_AND_M63_U1_nonlinearInst_n61), .A2(Fresh[33]), .ZN(
        top_AND_M63_U1_nonlinearInst_n62) );
  AND2_X1 top_AND_M63_U1_nonlinearInst_U22 ( .A1(Fresh[33]), .A2(
        top_AND_M63_U1_nonlinearInst_n61), .ZN(
        top_AND_M63_U1_nonlinearInst_n64) );
  OR2_X1 top_AND_M63_U1_nonlinearInst_U21 ( .A1(top_M41), .A2(top_T2), .ZN(
        top_AND_M63_U1_nonlinearInst_n61) );
  INV_X1 top_AND_M63_U1_nonlinearInst_U20 ( .A(top_AND_M63_U1_t[2]), .ZN(
        top_AND_M63_U1_t[6]) );
  OR2_X1 top_AND_M63_U1_nonlinearInst_U19 ( .A1(
        top_AND_M63_U1_nonlinearInst_n60), .A2(
        top_AND_M63_U1_nonlinearInst_n59), .ZN(top_AND_M63_U1_t[2]) );
  INV_X1 top_AND_M63_U1_nonlinearInst_U18 ( .A(
        top_AND_M63_U1_nonlinearInst_n58), .ZN(
        top_AND_M63_U1_nonlinearInst_n59) );
  OR2_X1 top_AND_M63_U1_nonlinearInst_U17 ( .A1(
        top_AND_M63_U1_nonlinearInst_n57), .A2(Fresh[33]), .ZN(
        top_AND_M63_U1_nonlinearInst_n58) );
  AND2_X1 top_AND_M63_U1_nonlinearInst_U16 ( .A1(Fresh[33]), .A2(
        top_AND_M63_U1_nonlinearInst_n57), .ZN(
        top_AND_M63_U1_nonlinearInst_n60) );
  OR2_X1 top_AND_M63_U1_nonlinearInst_U15 ( .A1(
        top_AND_M63_U1_nonlinearInst_n56), .A2(top_M41), .ZN(
        top_AND_M63_U1_nonlinearInst_n57) );
  INV_X1 top_AND_M63_U1_nonlinearInst_U14 ( .A(top_AND_M63_U1_t[1]), .ZN(
        top_AND_M63_U1_t[5]) );
  OR2_X1 top_AND_M63_U1_nonlinearInst_U13 ( .A1(
        top_AND_M63_U1_nonlinearInst_n55), .A2(
        top_AND_M63_U1_nonlinearInst_n54), .ZN(top_AND_M63_U1_t[1]) );
  AND2_X1 top_AND_M63_U1_nonlinearInst_U12 ( .A1(
        top_AND_M63_U1_nonlinearInst_n53), .A2(
        top_AND_M63_U1_nonlinearInst_n52), .ZN(
        top_AND_M63_U1_nonlinearInst_n54) );
  INV_X1 top_AND_M63_U1_nonlinearInst_U11 ( .A(
        top_AND_M63_U1_nonlinearInst_n51), .ZN(
        top_AND_M63_U1_nonlinearInst_n55) );
  OR2_X1 top_AND_M63_U1_nonlinearInst_U10 ( .A1(
        top_AND_M63_U1_nonlinearInst_n52), .A2(
        top_AND_M63_U1_nonlinearInst_n53), .ZN(
        top_AND_M63_U1_nonlinearInst_n51) );
  AND2_X1 top_AND_M63_U1_nonlinearInst_U9 ( .A1(top_M41), .A2(
        top_AND_M63_U1_nonlinearInst_n56), .ZN(
        top_AND_M63_U1_nonlinearInst_n53) );
  INV_X1 top_AND_M63_U1_nonlinearInst_U8 ( .A(top_T2), .ZN(
        top_AND_M63_U1_nonlinearInst_n56) );
  INV_X1 top_AND_M63_U1_nonlinearInst_U7 ( .A(top_AND_M63_U1_t[0]), .ZN(
        top_AND_M63_U1_t[4]) );
  OR2_X1 top_AND_M63_U1_nonlinearInst_U6 ( .A1(
        top_AND_M63_U1_nonlinearInst_n50), .A2(
        top_AND_M63_U1_nonlinearInst_n49), .ZN(top_AND_M63_U1_t[0]) );
  AND2_X1 top_AND_M63_U1_nonlinearInst_U5 ( .A1(
        top_AND_M63_U1_nonlinearInst_n48), .A2(
        top_AND_M63_U1_nonlinearInst_n52), .ZN(
        top_AND_M63_U1_nonlinearInst_n49) );
  INV_X1 top_AND_M63_U1_nonlinearInst_U4 ( .A(top_AND_M63_U1_nonlinearInst_n47), .ZN(top_AND_M63_U1_nonlinearInst_n50) );
  OR2_X1 top_AND_M63_U1_nonlinearInst_U3 ( .A1(
        top_AND_M63_U1_nonlinearInst_n52), .A2(
        top_AND_M63_U1_nonlinearInst_n48), .ZN(
        top_AND_M63_U1_nonlinearInst_n47) );
  AND2_X1 top_AND_M63_U1_nonlinearInst_U2 ( .A1(top_M41), .A2(top_T2), .ZN(
        top_AND_M63_U1_nonlinearInst_n48) );
  INV_X1 top_AND_M63_U1_nonlinearInst_U1 ( .A(Fresh[33]), .ZN(
        top_AND_M63_U1_nonlinearInst_n52) );
  AND2_X1 top_AND_M63_U1_gen_reg_0__regIns_U4 ( .A1(top_AND_M63_U1_t[0]), .A2(
        top_AND_M63_U1_gen_reg_0__regIns_n2), .ZN(
        top_AND_M63_U1_gen_reg_0__regIns_N3) );
  INV_X1 top_AND_M63_U1_gen_reg_0__regIns_U3 ( .A(reset), .ZN(
        top_AND_M63_U1_gen_reg_0__regIns_n2) );
  DFF_X1 top_AND_M63_U1_gen_reg_0__regIns_Q_reg ( .D(
        top_AND_M63_U1_gen_reg_0__regIns_N3), .CK(clk), .Q(
        top_AND_M63_U1_t_reg[0]) );
  AND2_X1 top_AND_M63_U1_gen_reg_1__regIns_U4 ( .A1(top_AND_M63_U1_t[1]), .A2(
        top_AND_M63_U1_gen_reg_1__regIns_n2), .ZN(
        top_AND_M63_U1_gen_reg_1__regIns_N3) );
  INV_X1 top_AND_M63_U1_gen_reg_1__regIns_U3 ( .A(reset), .ZN(
        top_AND_M63_U1_gen_reg_1__regIns_n2) );
  DFF_X1 top_AND_M63_U1_gen_reg_1__regIns_Q_reg ( .D(
        top_AND_M63_U1_gen_reg_1__regIns_N3), .CK(clk), .Q(
        top_AND_M63_U1_t_reg[1]) );
  AND2_X1 top_AND_M63_U1_gen_reg_2__regIns_U4 ( .A1(top_AND_M63_U1_t[2]), .A2(
        top_AND_M63_U1_gen_reg_2__regIns_n2), .ZN(
        top_AND_M63_U1_gen_reg_2__regIns_N3) );
  INV_X1 top_AND_M63_U1_gen_reg_2__regIns_U3 ( .A(reset), .ZN(
        top_AND_M63_U1_gen_reg_2__regIns_n2) );
  DFF_X1 top_AND_M63_U1_gen_reg_2__regIns_Q_reg ( .D(
        top_AND_M63_U1_gen_reg_2__regIns_N3), .CK(clk), .Q(
        top_AND_M63_U1_t_reg[2]) );
  AND2_X1 top_AND_M63_U1_gen_reg_3__regIns_U4 ( .A1(top_AND_M63_U1_t[3]), .A2(
        top_AND_M63_U1_gen_reg_3__regIns_n2), .ZN(
        top_AND_M63_U1_gen_reg_3__regIns_N3) );
  INV_X1 top_AND_M63_U1_gen_reg_3__regIns_U3 ( .A(reset), .ZN(
        top_AND_M63_U1_gen_reg_3__regIns_n2) );
  DFF_X1 top_AND_M63_U1_gen_reg_3__regIns_Q_reg ( .D(
        top_AND_M63_U1_gen_reg_3__regIns_N3), .CK(clk), .Q(
        top_AND_M63_U1_t_reg[3]) );
  AND2_X1 top_AND_M63_U1_gen_reg_4__regIns_U4 ( .A1(top_AND_M63_U1_t[4]), .A2(
        top_AND_M63_U1_gen_reg_4__regIns_n2), .ZN(
        top_AND_M63_U1_gen_reg_4__regIns_N3) );
  INV_X1 top_AND_M63_U1_gen_reg_4__regIns_U3 ( .A(reset), .ZN(
        top_AND_M63_U1_gen_reg_4__regIns_n2) );
  DFF_X1 top_AND_M63_U1_gen_reg_4__regIns_Q_reg ( .D(
        top_AND_M63_U1_gen_reg_4__regIns_N3), .CK(clk), .Q(
        top_AND_M63_U1_t_reg[4]) );
  AND2_X1 top_AND_M63_U1_gen_reg_5__regIns_U4 ( .A1(top_AND_M63_U1_t[5]), .A2(
        top_AND_M63_U1_gen_reg_5__regIns_n2), .ZN(
        top_AND_M63_U1_gen_reg_5__regIns_N3) );
  INV_X1 top_AND_M63_U1_gen_reg_5__regIns_U3 ( .A(reset), .ZN(
        top_AND_M63_U1_gen_reg_5__regIns_n2) );
  DFF_X1 top_AND_M63_U1_gen_reg_5__regIns_Q_reg ( .D(
        top_AND_M63_U1_gen_reg_5__regIns_N3), .CK(clk), .Q(
        top_AND_M63_U1_t_reg[5]) );
  AND2_X1 top_AND_M63_U1_gen_reg_6__regIns_U4 ( .A1(top_AND_M63_U1_t[6]), .A2(
        top_AND_M63_U1_gen_reg_6__regIns_n2), .ZN(
        top_AND_M63_U1_gen_reg_6__regIns_N3) );
  INV_X1 top_AND_M63_U1_gen_reg_6__regIns_U3 ( .A(reset), .ZN(
        top_AND_M63_U1_gen_reg_6__regIns_n2) );
  DFF_X1 top_AND_M63_U1_gen_reg_6__regIns_Q_reg ( .D(
        top_AND_M63_U1_gen_reg_6__regIns_N3), .CK(clk), .Q(
        top_AND_M63_U1_t_reg[6]) );
  AND2_X1 top_AND_M63_U1_gen_reg_7__regIns_U4 ( .A1(top_AND_M63_U1_t[7]), .A2(
        top_AND_M63_U1_gen_reg_7__regIns_n2), .ZN(
        top_AND_M63_U1_gen_reg_7__regIns_N3) );
  INV_X1 top_AND_M63_U1_gen_reg_7__regIns_U3 ( .A(reset), .ZN(
        top_AND_M63_U1_gen_reg_7__regIns_n2) );
  DFF_X1 top_AND_M63_U1_gen_reg_7__regIns_Q_reg ( .D(
        top_AND_M63_U1_gen_reg_7__regIns_N3), .CK(clk), .Q(
        top_AND_M63_U1_t_reg[7]) );
  AND2_X1 top_AND_M63_U1_OperationInst_andInst0_U2 ( .A1(
        top_new_AGEMA_signal_164), .A2(
        top_AND_M63_U1_OperationInst_andInst0_n3), .ZN(
        top_AND_M63_U1_OperationInst_q[0]) );
  AND2_X1 top_AND_M63_U1_OperationInst_andInst0_U1 ( .A1(
        top_new_AGEMA_signal_306), .A2(top_AND_M63_U1_t_reg[0]), .ZN(
        top_AND_M63_U1_OperationInst_andInst0_n3) );
  AND2_X1 top_AND_M63_U1_OperationInst_andInst1_U2 ( .A1(
        top_new_AGEMA_signal_163), .A2(
        top_AND_M63_U1_OperationInst_andInst1_n3), .ZN(
        top_AND_M63_U1_OperationInst_q[1]) );
  AND2_X1 top_AND_M63_U1_OperationInst_andInst1_U1 ( .A1(
        top_new_AGEMA_signal_306), .A2(top_AND_M63_U1_t_reg[1]), .ZN(
        top_AND_M63_U1_OperationInst_andInst1_n3) );
  AND2_X1 top_AND_M63_U1_OperationInst_andInst2_U2 ( .A1(
        top_new_AGEMA_signal_164), .A2(
        top_AND_M63_U1_OperationInst_andInst2_n3), .ZN(
        top_AND_M63_U1_OperationInst_q[2]) );
  AND2_X1 top_AND_M63_U1_OperationInst_andInst2_U1 ( .A1(
        top_new_AGEMA_signal_305), .A2(top_AND_M63_U1_t_reg[2]), .ZN(
        top_AND_M63_U1_OperationInst_andInst2_n3) );
  AND2_X1 top_AND_M63_U1_OperationInst_andInst3_U2 ( .A1(
        top_new_AGEMA_signal_163), .A2(
        top_AND_M63_U1_OperationInst_andInst3_n3), .ZN(
        top_AND_M63_U1_OperationInst_q[3]) );
  AND2_X1 top_AND_M63_U1_OperationInst_andInst3_U1 ( .A1(
        top_new_AGEMA_signal_305), .A2(top_AND_M63_U1_t_reg[3]), .ZN(
        top_AND_M63_U1_OperationInst_andInst3_n3) );
  OR2_X1 top_AND_M63_U1_OperationInst_orInst1_U3 ( .A1(
        top_AND_M63_U1_OperationInst_q[1]), .A2(
        top_AND_M63_U1_OperationInst_orInst1_n6), .ZN(top_new_AGEMA_signal_345) );
  OR2_X1 top_AND_M63_U1_OperationInst_orInst1_U2 ( .A1(
        top_AND_M63_U1_OperationInst_q[0]), .A2(
        top_AND_M63_U1_OperationInst_orInst1_n5), .ZN(
        top_AND_M63_U1_OperationInst_orInst1_n6) );
  OR2_X1 top_AND_M63_U1_OperationInst_orInst1_U1 ( .A1(
        top_AND_M63_U1_OperationInst_q[3]), .A2(
        top_AND_M63_U1_OperationInst_q[2]), .ZN(
        top_AND_M63_U1_OperationInst_orInst1_n5) );
  AND2_X1 top_AND_M63_U1_OperationInst_andInst4_U2 ( .A1(
        top_new_AGEMA_signal_164), .A2(
        top_AND_M63_U1_OperationInst_andInst4_n3), .ZN(
        top_AND_M63_U1_OperationInst_q[4]) );
  AND2_X1 top_AND_M63_U1_OperationInst_andInst4_U1 ( .A1(
        top_new_AGEMA_signal_306), .A2(top_AND_M63_U1_t_reg[4]), .ZN(
        top_AND_M63_U1_OperationInst_andInst4_n3) );
  AND2_X1 top_AND_M63_U1_OperationInst_andInst5_U2 ( .A1(
        top_new_AGEMA_signal_163), .A2(
        top_AND_M63_U1_OperationInst_andInst5_n3), .ZN(
        top_AND_M63_U1_OperationInst_q[5]) );
  AND2_X1 top_AND_M63_U1_OperationInst_andInst5_U1 ( .A1(
        top_new_AGEMA_signal_306), .A2(top_AND_M63_U1_t_reg[5]), .ZN(
        top_AND_M63_U1_OperationInst_andInst5_n3) );
  AND2_X1 top_AND_M63_U1_OperationInst_andInst6_U2 ( .A1(
        top_new_AGEMA_signal_164), .A2(
        top_AND_M63_U1_OperationInst_andInst6_n3), .ZN(
        top_AND_M63_U1_OperationInst_q[6]) );
  AND2_X1 top_AND_M63_U1_OperationInst_andInst6_U1 ( .A1(
        top_new_AGEMA_signal_305), .A2(top_AND_M63_U1_t_reg[6]), .ZN(
        top_AND_M63_U1_OperationInst_andInst6_n3) );
  AND2_X1 top_AND_M63_U1_OperationInst_andInst7_U2 ( .A1(
        top_new_AGEMA_signal_163), .A2(
        top_AND_M63_U1_OperationInst_andInst7_n3), .ZN(
        top_AND_M63_U1_OperationInst_q[7]) );
  AND2_X1 top_AND_M63_U1_OperationInst_andInst7_U1 ( .A1(
        top_new_AGEMA_signal_305), .A2(top_AND_M63_U1_t_reg[7]), .ZN(
        top_AND_M63_U1_OperationInst_andInst7_n3) );
  OR2_X1 top_AND_M63_U1_OperationInst_orInst2_U3 ( .A1(
        top_AND_M63_U1_OperationInst_q[5]), .A2(
        top_AND_M63_U1_OperationInst_orInst2_n6), .ZN(top_new_AGEMA_signal_346) );
  OR2_X1 top_AND_M63_U1_OperationInst_orInst2_U2 ( .A1(
        top_AND_M63_U1_OperationInst_q[4]), .A2(
        top_AND_M63_U1_OperationInst_orInst2_n5), .ZN(
        top_AND_M63_U1_OperationInst_orInst2_n6) );
  OR2_X1 top_AND_M63_U1_OperationInst_orInst2_U1 ( .A1(
        top_AND_M63_U1_OperationInst_q[7]), .A2(
        top_AND_M63_U1_OperationInst_q[6]), .ZN(
        top_AND_M63_U1_OperationInst_orInst2_n5) );
  OR2_X1 top_XOR_L0_U1_xorInst_U5 ( .A1(top_XOR_L0_U1_xorInst_n12), .A2(
        top_XOR_L0_U1_xorInst_n11), .ZN(top_L0) );
  INV_X1 top_XOR_L0_U1_xorInst_U4 ( .A(top_XOR_L0_U1_xorInst_n10), .ZN(
        top_XOR_L0_U1_xorInst_n11) );
  OR2_X1 top_XOR_L0_U1_xorInst_U3 ( .A1(top_XOR_L0_U1_xorInst_n9), .A2(
        Fresh[31]), .ZN(top_XOR_L0_U1_xorInst_n10) );
  AND2_X1 top_XOR_L0_U1_xorInst_U2 ( .A1(Fresh[31]), .A2(
        top_XOR_L0_U1_xorInst_n9), .ZN(top_XOR_L0_U1_xorInst_n12) );
  INV_X1 top_XOR_L0_U1_xorInst_U1 ( .A(Fresh[32]), .ZN(
        top_XOR_L0_U1_xorInst_n9) );
  AND2_X1 top_XOR_L0_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_355), .A2(
        top_new_AGEMA_signal_344), .ZN(top_XOR_L0_U1_w[0]) );
  AND2_X1 top_XOR_L0_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_356), .A2(
        top_new_AGEMA_signal_343), .ZN(top_XOR_L0_U1_w[1]) );
  AND2_X1 top_XOR_L0_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_356), .A2(
        top_new_AGEMA_signal_344), .ZN(top_XOR_L0_U1_w[2]) );
  AND2_X1 top_XOR_L0_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_355), .A2(
        top_new_AGEMA_signal_343), .ZN(top_XOR_L0_U1_w[3]) );
  OR2_X1 top_XOR_L0_U1_orInst1_U1 ( .A1(top_XOR_L0_U1_w[0]), .A2(
        top_XOR_L0_U1_w[1]), .ZN(top_new_AGEMA_signal_373) );
  OR2_X1 top_XOR_L0_U1_orInst2_U1 ( .A1(top_XOR_L0_U1_w[2]), .A2(
        top_XOR_L0_U1_w[3]), .ZN(top_new_AGEMA_signal_374) );
  OR2_X1 top_XOR_L1_U1_xorInst_U5 ( .A1(top_XOR_L1_U1_xorInst_n12), .A2(
        top_XOR_L1_U1_xorInst_n11), .ZN(top_L1) );
  INV_X1 top_XOR_L1_U1_xorInst_U4 ( .A(top_XOR_L1_U1_xorInst_n10), .ZN(
        top_XOR_L1_U1_xorInst_n11) );
  OR2_X1 top_XOR_L1_U1_xorInst_U3 ( .A1(top_XOR_L1_U1_xorInst_n9), .A2(
        Fresh[20]), .ZN(top_XOR_L1_U1_xorInst_n10) );
  AND2_X1 top_XOR_L1_U1_xorInst_U2 ( .A1(Fresh[20]), .A2(
        top_XOR_L1_U1_xorInst_n9), .ZN(top_XOR_L1_U1_xorInst_n12) );
  INV_X1 top_XOR_L1_U1_xorInst_U1 ( .A(Fresh[26]), .ZN(
        top_XOR_L1_U1_xorInst_n9) );
  AND2_X1 top_XOR_L1_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_321), .A2(
        top_new_AGEMA_signal_318), .ZN(top_XOR_L1_U1_w[0]) );
  AND2_X1 top_XOR_L1_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_322), .A2(
        top_new_AGEMA_signal_317), .ZN(top_XOR_L1_U1_w[1]) );
  AND2_X1 top_XOR_L1_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_322), .A2(
        top_new_AGEMA_signal_318), .ZN(top_XOR_L1_U1_w[2]) );
  AND2_X1 top_XOR_L1_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_321), .A2(
        top_new_AGEMA_signal_317), .ZN(top_XOR_L1_U1_w[3]) );
  OR2_X1 top_XOR_L1_U1_orInst1_U1 ( .A1(top_XOR_L1_U1_w[0]), .A2(
        top_XOR_L1_U1_w[1]), .ZN(top_new_AGEMA_signal_347) );
  OR2_X1 top_XOR_L1_U1_orInst2_U1 ( .A1(top_XOR_L1_U1_w[2]), .A2(
        top_XOR_L1_U1_w[3]), .ZN(top_new_AGEMA_signal_348) );
  OR2_X1 top_XOR_L2_U1_xorInst_U5 ( .A1(top_XOR_L2_U1_xorInst_n12), .A2(
        top_XOR_L2_U1_xorInst_n11), .ZN(top_L2) );
  INV_X1 top_XOR_L2_U1_xorInst_U4 ( .A(top_XOR_L2_U1_xorInst_n10), .ZN(
        top_XOR_L2_U1_xorInst_n11) );
  OR2_X1 top_XOR_L2_U1_xorInst_U3 ( .A1(top_XOR_L2_U1_xorInst_n9), .A2(
        Fresh[16]), .ZN(top_XOR_L2_U1_xorInst_n10) );
  AND2_X1 top_XOR_L2_U1_xorInst_U2 ( .A1(Fresh[16]), .A2(
        top_XOR_L2_U1_xorInst_n9), .ZN(top_XOR_L2_U1_xorInst_n12) );
  INV_X1 top_XOR_L2_U1_xorInst_U1 ( .A(Fresh[18]), .ZN(
        top_XOR_L2_U1_xorInst_n9) );
  AND2_X1 top_XOR_L2_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_315), .A2(
        top_new_AGEMA_signal_332), .ZN(top_XOR_L2_U1_w[0]) );
  AND2_X1 top_XOR_L2_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_316), .A2(
        top_new_AGEMA_signal_331), .ZN(top_XOR_L2_U1_w[1]) );
  AND2_X1 top_XOR_L2_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_316), .A2(
        top_new_AGEMA_signal_332), .ZN(top_XOR_L2_U1_w[2]) );
  AND2_X1 top_XOR_L2_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_315), .A2(
        top_new_AGEMA_signal_331), .ZN(top_XOR_L2_U1_w[3]) );
  OR2_X1 top_XOR_L2_U1_orInst1_U1 ( .A1(top_XOR_L2_U1_w[0]), .A2(
        top_XOR_L2_U1_w[1]), .ZN(top_new_AGEMA_signal_357) );
  OR2_X1 top_XOR_L2_U1_orInst2_U1 ( .A1(top_XOR_L2_U1_w[2]), .A2(
        top_XOR_L2_U1_w[3]), .ZN(top_new_AGEMA_signal_358) );
  OR2_X1 top_XOR_L3_U1_xorInst_U5 ( .A1(top_XOR_L3_U1_xorInst_n12), .A2(
        top_XOR_L3_U1_xorInst_n11), .ZN(top_L3) );
  INV_X1 top_XOR_L3_U1_xorInst_U4 ( .A(top_XOR_L3_U1_xorInst_n10), .ZN(
        top_XOR_L3_U1_xorInst_n11) );
  OR2_X1 top_XOR_L3_U1_xorInst_U3 ( .A1(top_XOR_L3_U1_xorInst_n9), .A2(
        Fresh[17]), .ZN(top_XOR_L3_U1_xorInst_n10) );
  AND2_X1 top_XOR_L3_U1_xorInst_U2 ( .A1(Fresh[17]), .A2(
        top_XOR_L3_U1_xorInst_n9), .ZN(top_XOR_L3_U1_xorInst_n12) );
  INV_X1 top_XOR_L3_U1_xorInst_U1 ( .A(Fresh[25]), .ZN(
        top_XOR_L3_U1_xorInst_n9) );
  AND2_X1 top_XOR_L3_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_339), .A2(
        top_new_AGEMA_signal_314), .ZN(top_XOR_L3_U1_w[0]) );
  AND2_X1 top_XOR_L3_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_340), .A2(
        top_new_AGEMA_signal_313), .ZN(top_XOR_L3_U1_w[1]) );
  AND2_X1 top_XOR_L3_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_340), .A2(
        top_new_AGEMA_signal_314), .ZN(top_XOR_L3_U1_w[2]) );
  AND2_X1 top_XOR_L3_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_339), .A2(
        top_new_AGEMA_signal_313), .ZN(top_XOR_L3_U1_w[3]) );
  OR2_X1 top_XOR_L3_U1_orInst1_U1 ( .A1(top_XOR_L3_U1_w[0]), .A2(
        top_XOR_L3_U1_w[1]), .ZN(top_new_AGEMA_signal_359) );
  OR2_X1 top_XOR_L3_U1_orInst2_U1 ( .A1(top_XOR_L3_U1_w[2]), .A2(
        top_XOR_L3_U1_w[3]), .ZN(top_new_AGEMA_signal_360) );
  OR2_X1 top_XOR_L4_U1_xorInst_U5 ( .A1(top_XOR_L4_U1_xorInst_n12), .A2(
        top_XOR_L4_U1_xorInst_n11), .ZN(top_L4) );
  INV_X1 top_XOR_L4_U1_xorInst_U4 ( .A(top_XOR_L4_U1_xorInst_n10), .ZN(
        top_XOR_L4_U1_xorInst_n11) );
  OR2_X1 top_XOR_L4_U1_xorInst_U3 ( .A1(top_XOR_L4_U1_xorInst_n9), .A2(
        Fresh[24]), .ZN(top_XOR_L4_U1_xorInst_n10) );
  AND2_X1 top_XOR_L4_U1_xorInst_U2 ( .A1(Fresh[24]), .A2(
        top_XOR_L4_U1_xorInst_n9), .ZN(top_XOR_L4_U1_xorInst_n12) );
  INV_X1 top_XOR_L4_U1_xorInst_U1 ( .A(Fresh[28]), .ZN(
        top_XOR_L4_U1_xorInst_n9) );
  AND2_X1 top_XOR_L4_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_341), .A2(
        top_new_AGEMA_signal_338), .ZN(top_XOR_L4_U1_w[0]) );
  AND2_X1 top_XOR_L4_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_342), .A2(
        top_new_AGEMA_signal_337), .ZN(top_XOR_L4_U1_w[1]) );
  AND2_X1 top_XOR_L4_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_342), .A2(
        top_new_AGEMA_signal_338), .ZN(top_XOR_L4_U1_w[2]) );
  AND2_X1 top_XOR_L4_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_341), .A2(
        top_new_AGEMA_signal_337), .ZN(top_XOR_L4_U1_w[3]) );
  OR2_X1 top_XOR_L4_U1_orInst1_U1 ( .A1(top_XOR_L4_U1_w[0]), .A2(
        top_XOR_L4_U1_w[1]), .ZN(top_new_AGEMA_signal_361) );
  OR2_X1 top_XOR_L4_U1_orInst2_U1 ( .A1(top_XOR_L4_U1_w[2]), .A2(
        top_XOR_L4_U1_w[3]), .ZN(top_new_AGEMA_signal_362) );
  OR2_X1 top_XOR_L5_U1_xorInst_U5 ( .A1(top_XOR_L5_U1_xorInst_n12), .A2(
        top_XOR_L5_U1_xorInst_n11), .ZN(top_L5) );
  INV_X1 top_XOR_L5_U1_xorInst_U4 ( .A(top_XOR_L5_U1_xorInst_n10), .ZN(
        top_XOR_L5_U1_xorInst_n11) );
  OR2_X1 top_XOR_L5_U1_xorInst_U3 ( .A1(top_XOR_L5_U1_xorInst_n9), .A2(
        Fresh[19]), .ZN(top_XOR_L5_U1_xorInst_n10) );
  AND2_X1 top_XOR_L5_U1_xorInst_U2 ( .A1(Fresh[19]), .A2(
        top_XOR_L5_U1_xorInst_n9), .ZN(top_XOR_L5_U1_xorInst_n12) );
  INV_X1 top_XOR_L5_U1_xorInst_U1 ( .A(Fresh[31]), .ZN(
        top_XOR_L5_U1_xorInst_n9) );
  AND2_X1 top_XOR_L5_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_343), .A2(
        top_new_AGEMA_signal_334), .ZN(top_XOR_L5_U1_w[0]) );
  AND2_X1 top_XOR_L5_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_344), .A2(
        top_new_AGEMA_signal_333), .ZN(top_XOR_L5_U1_w[1]) );
  AND2_X1 top_XOR_L5_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_344), .A2(
        top_new_AGEMA_signal_334), .ZN(top_XOR_L5_U1_w[2]) );
  AND2_X1 top_XOR_L5_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_343), .A2(
        top_new_AGEMA_signal_333), .ZN(top_XOR_L5_U1_w[3]) );
  OR2_X1 top_XOR_L5_U1_orInst1_U1 ( .A1(top_XOR_L5_U1_w[0]), .A2(
        top_XOR_L5_U1_w[1]), .ZN(top_new_AGEMA_signal_363) );
  OR2_X1 top_XOR_L5_U1_orInst2_U1 ( .A1(top_XOR_L5_U1_w[2]), .A2(
        top_XOR_L5_U1_w[3]), .ZN(top_new_AGEMA_signal_364) );
  OR2_X1 top_XOR_L6_U1_xorInst_U5 ( .A1(top_XOR_L6_U1_xorInst_n12), .A2(
        top_XOR_L6_U1_xorInst_n11), .ZN(top_L6) );
  INV_X1 top_XOR_L6_U1_xorInst_U4 ( .A(top_XOR_L6_U1_xorInst_n10), .ZN(
        top_XOR_L6_U1_xorInst_n11) );
  OR2_X1 top_XOR_L6_U1_xorInst_U3 ( .A1(top_XOR_L6_U1_xorInst_n9), .A2(
        Fresh[32]), .ZN(top_XOR_L6_U1_xorInst_n10) );
  AND2_X1 top_XOR_L6_U1_xorInst_U2 ( .A1(Fresh[32]), .A2(
        top_XOR_L6_U1_xorInst_n9), .ZN(top_XOR_L6_U1_xorInst_n12) );
  INV_X1 top_XOR_L6_U1_xorInst_U1 ( .A(top_L5), .ZN(top_XOR_L6_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_L6_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_363), .A2(
        top_new_AGEMA_signal_356), .ZN(top_XOR_L6_U1_w[0]) );
  AND2_X1 top_XOR_L6_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_364), .A2(
        top_new_AGEMA_signal_355), .ZN(top_XOR_L6_U1_w[1]) );
  AND2_X1 top_XOR_L6_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_364), .A2(
        top_new_AGEMA_signal_356), .ZN(top_XOR_L6_U1_w[2]) );
  AND2_X1 top_XOR_L6_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_363), .A2(
        top_new_AGEMA_signal_355), .ZN(top_XOR_L6_U1_w[3]) );
  OR2_X1 top_XOR_L6_U1_orInst1_U1 ( .A1(top_XOR_L6_U1_w[0]), .A2(
        top_XOR_L6_U1_w[1]), .ZN(top_new_AGEMA_signal_375) );
  OR2_X1 top_XOR_L6_U1_orInst2_U1 ( .A1(top_XOR_L6_U1_w[2]), .A2(
        top_XOR_L6_U1_w[3]), .ZN(top_new_AGEMA_signal_376) );
  OR2_X1 top_XOR_L7_U1_xorInst_U5 ( .A1(top_XOR_L7_U1_xorInst_n12), .A2(
        top_XOR_L7_U1_xorInst_n11), .ZN(top_L7) );
  INV_X1 top_XOR_L7_U1_xorInst_U4 ( .A(top_XOR_L7_U1_xorInst_n10), .ZN(
        top_XOR_L7_U1_xorInst_n11) );
  OR2_X1 top_XOR_L7_U1_xorInst_U3 ( .A1(top_XOR_L7_U1_xorInst_n9), .A2(
        Fresh[16]), .ZN(top_XOR_L7_U1_xorInst_n10) );
  AND2_X1 top_XOR_L7_U1_xorInst_U2 ( .A1(Fresh[16]), .A2(
        top_XOR_L7_U1_xorInst_n9), .ZN(top_XOR_L7_U1_xorInst_n12) );
  INV_X1 top_XOR_L7_U1_xorInst_U1 ( .A(top_L3), .ZN(top_XOR_L7_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_L7_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_359), .A2(
        top_new_AGEMA_signal_332), .ZN(top_XOR_L7_U1_w[0]) );
  AND2_X1 top_XOR_L7_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_360), .A2(
        top_new_AGEMA_signal_331), .ZN(top_XOR_L7_U1_w[1]) );
  AND2_X1 top_XOR_L7_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_360), .A2(
        top_new_AGEMA_signal_332), .ZN(top_XOR_L7_U1_w[2]) );
  AND2_X1 top_XOR_L7_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_359), .A2(
        top_new_AGEMA_signal_331), .ZN(top_XOR_L7_U1_w[3]) );
  OR2_X1 top_XOR_L7_U1_orInst1_U1 ( .A1(top_XOR_L7_U1_w[0]), .A2(
        top_XOR_L7_U1_w[1]), .ZN(top_new_AGEMA_signal_377) );
  OR2_X1 top_XOR_L7_U1_orInst2_U1 ( .A1(top_XOR_L7_U1_w[2]), .A2(
        top_XOR_L7_U1_w[3]), .ZN(top_new_AGEMA_signal_378) );
  OR2_X1 top_XOR_L8_U1_xorInst_U5 ( .A1(top_XOR_L8_U1_xorInst_n12), .A2(
        top_XOR_L8_U1_xorInst_n11), .ZN(top_L8) );
  INV_X1 top_XOR_L8_U1_xorInst_U4 ( .A(top_XOR_L8_U1_xorInst_n10), .ZN(
        top_XOR_L8_U1_xorInst_n11) );
  OR2_X1 top_XOR_L8_U1_xorInst_U3 ( .A1(top_XOR_L8_U1_xorInst_n9), .A2(
        Fresh[21]), .ZN(top_XOR_L8_U1_xorInst_n10) );
  AND2_X1 top_XOR_L8_U1_xorInst_U2 ( .A1(Fresh[21]), .A2(
        top_XOR_L8_U1_xorInst_n9), .ZN(top_XOR_L8_U1_xorInst_n12) );
  INV_X1 top_XOR_L8_U1_xorInst_U1 ( .A(Fresh[29]), .ZN(
        top_XOR_L8_U1_xorInst_n9) );
  AND2_X1 top_XOR_L8_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_325), .A2(
        top_new_AGEMA_signal_320), .ZN(top_XOR_L8_U1_w[0]) );
  AND2_X1 top_XOR_L8_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_326), .A2(
        top_new_AGEMA_signal_319), .ZN(top_XOR_L8_U1_w[1]) );
  AND2_X1 top_XOR_L8_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_326), .A2(
        top_new_AGEMA_signal_320), .ZN(top_XOR_L8_U1_w[2]) );
  AND2_X1 top_XOR_L8_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_325), .A2(
        top_new_AGEMA_signal_319), .ZN(top_XOR_L8_U1_w[3]) );
  OR2_X1 top_XOR_L8_U1_orInst1_U1 ( .A1(top_XOR_L8_U1_w[0]), .A2(
        top_XOR_L8_U1_w[1]), .ZN(top_new_AGEMA_signal_349) );
  OR2_X1 top_XOR_L8_U1_orInst2_U1 ( .A1(top_XOR_L8_U1_w[2]), .A2(
        top_XOR_L8_U1_w[3]), .ZN(top_new_AGEMA_signal_350) );
  OR2_X1 top_XOR_L9_U1_xorInst_U5 ( .A1(top_XOR_L9_U1_xorInst_n12), .A2(
        top_XOR_L9_U1_xorInst_n11), .ZN(top_L9) );
  INV_X1 top_XOR_L9_U1_xorInst_U4 ( .A(top_XOR_L9_U1_xorInst_n10), .ZN(
        top_XOR_L9_U1_xorInst_n11) );
  OR2_X1 top_XOR_L9_U1_xorInst_U3 ( .A1(top_XOR_L9_U1_xorInst_n9), .A2(
        Fresh[22]), .ZN(top_XOR_L9_U1_xorInst_n10) );
  AND2_X1 top_XOR_L9_U1_xorInst_U2 ( .A1(Fresh[22]), .A2(
        top_XOR_L9_U1_xorInst_n9), .ZN(top_XOR_L9_U1_xorInst_n12) );
  INV_X1 top_XOR_L9_U1_xorInst_U1 ( .A(Fresh[23]), .ZN(
        top_XOR_L9_U1_xorInst_n9) );
  AND2_X1 top_XOR_L9_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_353), .A2(
        top_new_AGEMA_signal_336), .ZN(top_XOR_L9_U1_w[0]) );
  AND2_X1 top_XOR_L9_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_354), .A2(
        top_new_AGEMA_signal_335), .ZN(top_XOR_L9_U1_w[1]) );
  AND2_X1 top_XOR_L9_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_354), .A2(
        top_new_AGEMA_signal_336), .ZN(top_XOR_L9_U1_w[2]) );
  AND2_X1 top_XOR_L9_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_353), .A2(
        top_new_AGEMA_signal_335), .ZN(top_XOR_L9_U1_w[3]) );
  OR2_X1 top_XOR_L9_U1_orInst1_U1 ( .A1(top_XOR_L9_U1_w[0]), .A2(
        top_XOR_L9_U1_w[1]), .ZN(top_new_AGEMA_signal_379) );
  OR2_X1 top_XOR_L9_U1_orInst2_U1 ( .A1(top_XOR_L9_U1_w[2]), .A2(
        top_XOR_L9_U1_w[3]), .ZN(top_new_AGEMA_signal_380) );
  OR2_X1 top_XOR_L10_U1_xorInst_U5 ( .A1(top_XOR_L10_U1_xorInst_n12), .A2(
        top_XOR_L10_U1_xorInst_n11), .ZN(top_L10) );
  INV_X1 top_XOR_L10_U1_xorInst_U4 ( .A(top_XOR_L10_U1_xorInst_n10), .ZN(
        top_XOR_L10_U1_xorInst_n11) );
  OR2_X1 top_XOR_L10_U1_xorInst_U3 ( .A1(top_XOR_L10_U1_xorInst_n9), .A2(
        Fresh[23]), .ZN(top_XOR_L10_U1_xorInst_n10) );
  AND2_X1 top_XOR_L10_U1_xorInst_U2 ( .A1(Fresh[23]), .A2(
        top_XOR_L10_U1_xorInst_n9), .ZN(top_XOR_L10_U1_xorInst_n12) );
  INV_X1 top_XOR_L10_U1_xorInst_U1 ( .A(top_L4), .ZN(top_XOR_L10_U1_xorInst_n9) );
  AND2_X1 top_XOR_L10_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_361), .A2(
        top_new_AGEMA_signal_354), .ZN(top_XOR_L10_U1_w[0]) );
  AND2_X1 top_XOR_L10_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_362), .A2(
        top_new_AGEMA_signal_353), .ZN(top_XOR_L10_U1_w[1]) );
  AND2_X1 top_XOR_L10_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_362), .A2(
        top_new_AGEMA_signal_354), .ZN(top_XOR_L10_U1_w[2]) );
  AND2_X1 top_XOR_L10_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_361), .A2(
        top_new_AGEMA_signal_353), .ZN(top_XOR_L10_U1_w[3]) );
  OR2_X1 top_XOR_L10_U1_orInst1_U1 ( .A1(top_XOR_L10_U1_w[0]), .A2(
        top_XOR_L10_U1_w[1]), .ZN(top_new_AGEMA_signal_381) );
  OR2_X1 top_XOR_L10_U1_orInst2_U1 ( .A1(top_XOR_L10_U1_w[2]), .A2(
        top_XOR_L10_U1_w[3]), .ZN(top_new_AGEMA_signal_382) );
  OR2_X1 top_XOR_L11_U1_xorInst_U5 ( .A1(top_XOR_L11_U1_xorInst_n12), .A2(
        top_XOR_L11_U1_xorInst_n11), .ZN(top_L11) );
  INV_X1 top_XOR_L11_U1_xorInst_U4 ( .A(top_XOR_L11_U1_xorInst_n10), .ZN(
        top_XOR_L11_U1_xorInst_n11) );
  OR2_X1 top_XOR_L11_U1_xorInst_U3 ( .A1(top_XOR_L11_U1_xorInst_n9), .A2(
        Fresh[30]), .ZN(top_XOR_L11_U1_xorInst_n10) );
  AND2_X1 top_XOR_L11_U1_xorInst_U2 ( .A1(Fresh[30]), .A2(
        top_XOR_L11_U1_xorInst_n9), .ZN(top_XOR_L11_U1_xorInst_n12) );
  INV_X1 top_XOR_L11_U1_xorInst_U1 ( .A(top_L2), .ZN(top_XOR_L11_U1_xorInst_n9) );
  AND2_X1 top_XOR_L11_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_357), .A2(
        top_new_AGEMA_signal_328), .ZN(top_XOR_L11_U1_w[0]) );
  AND2_X1 top_XOR_L11_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_358), .A2(
        top_new_AGEMA_signal_327), .ZN(top_XOR_L11_U1_w[1]) );
  AND2_X1 top_XOR_L11_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_358), .A2(
        top_new_AGEMA_signal_328), .ZN(top_XOR_L11_U1_w[2]) );
  AND2_X1 top_XOR_L11_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_357), .A2(
        top_new_AGEMA_signal_327), .ZN(top_XOR_L11_U1_w[3]) );
  OR2_X1 top_XOR_L11_U1_orInst1_U1 ( .A1(top_XOR_L11_U1_w[0]), .A2(
        top_XOR_L11_U1_w[1]), .ZN(top_new_AGEMA_signal_383) );
  OR2_X1 top_XOR_L11_U1_orInst2_U1 ( .A1(top_XOR_L11_U1_w[2]), .A2(
        top_XOR_L11_U1_w[3]), .ZN(top_new_AGEMA_signal_384) );
  OR2_X1 top_XOR_L12_U1_xorInst_U5 ( .A1(top_XOR_L12_U1_xorInst_n12), .A2(
        top_XOR_L12_U1_xorInst_n11), .ZN(top_L12) );
  INV_X1 top_XOR_L12_U1_xorInst_U4 ( .A(top_XOR_L12_U1_xorInst_n10), .ZN(
        top_XOR_L12_U1_xorInst_n11) );
  OR2_X1 top_XOR_L12_U1_xorInst_U3 ( .A1(top_XOR_L12_U1_xorInst_n9), .A2(
        Fresh[18]), .ZN(top_XOR_L12_U1_xorInst_n10) );
  AND2_X1 top_XOR_L12_U1_xorInst_U2 ( .A1(Fresh[18]), .A2(
        top_XOR_L12_U1_xorInst_n9), .ZN(top_XOR_L12_U1_xorInst_n12) );
  INV_X1 top_XOR_L12_U1_xorInst_U1 ( .A(Fresh[21]), .ZN(
        top_XOR_L12_U1_xorInst_n9) );
  AND2_X1 top_XOR_L12_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_319), .A2(
        top_new_AGEMA_signal_316), .ZN(top_XOR_L12_U1_w[0]) );
  AND2_X1 top_XOR_L12_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_320), .A2(
        top_new_AGEMA_signal_315), .ZN(top_XOR_L12_U1_w[1]) );
  AND2_X1 top_XOR_L12_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_320), .A2(
        top_new_AGEMA_signal_316), .ZN(top_XOR_L12_U1_w[2]) );
  AND2_X1 top_XOR_L12_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_319), .A2(
        top_new_AGEMA_signal_315), .ZN(top_XOR_L12_U1_w[3]) );
  OR2_X1 top_XOR_L12_U1_orInst1_U1 ( .A1(top_XOR_L12_U1_w[0]), .A2(
        top_XOR_L12_U1_w[1]), .ZN(top_new_AGEMA_signal_351) );
  OR2_X1 top_XOR_L12_U1_orInst2_U1 ( .A1(top_XOR_L12_U1_w[2]), .A2(
        top_XOR_L12_U1_w[3]), .ZN(top_new_AGEMA_signal_352) );
  OR2_X1 top_XOR_L13_U1_xorInst_U5 ( .A1(top_XOR_L13_U1_xorInst_n12), .A2(
        top_XOR_L13_U1_xorInst_n11), .ZN(top_L13) );
  INV_X1 top_XOR_L13_U1_xorInst_U4 ( .A(top_XOR_L13_U1_xorInst_n10), .ZN(
        top_XOR_L13_U1_xorInst_n11) );
  OR2_X1 top_XOR_L13_U1_xorInst_U3 ( .A1(top_XOR_L13_U1_xorInst_n9), .A2(
        Fresh[20]), .ZN(top_XOR_L13_U1_xorInst_n10) );
  AND2_X1 top_XOR_L13_U1_xorInst_U2 ( .A1(Fresh[20]), .A2(
        top_XOR_L13_U1_xorInst_n9), .ZN(top_XOR_L13_U1_xorInst_n12) );
  INV_X1 top_XOR_L13_U1_xorInst_U1 ( .A(top_L0), .ZN(top_XOR_L13_U1_xorInst_n9) );
  AND2_X1 top_XOR_L13_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_373), .A2(
        top_new_AGEMA_signal_318), .ZN(top_XOR_L13_U1_w[0]) );
  AND2_X1 top_XOR_L13_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_374), .A2(
        top_new_AGEMA_signal_317), .ZN(top_XOR_L13_U1_w[1]) );
  AND2_X1 top_XOR_L13_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_374), .A2(
        top_new_AGEMA_signal_318), .ZN(top_XOR_L13_U1_w[2]) );
  AND2_X1 top_XOR_L13_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_373), .A2(
        top_new_AGEMA_signal_317), .ZN(top_XOR_L13_U1_w[3]) );
  OR2_X1 top_XOR_L13_U1_orInst1_U1 ( .A1(top_XOR_L13_U1_w[0]), .A2(
        top_XOR_L13_U1_w[1]), .ZN(top_new_AGEMA_signal_391) );
  OR2_X1 top_XOR_L13_U1_orInst2_U1 ( .A1(top_XOR_L13_U1_w[2]), .A2(
        top_XOR_L13_U1_w[3]), .ZN(top_new_AGEMA_signal_392) );
  OR2_X1 top_XOR_L14_U1_xorInst_U5 ( .A1(top_XOR_L14_U1_xorInst_n12), .A2(
        top_XOR_L14_U1_xorInst_n11), .ZN(top_L14) );
  INV_X1 top_XOR_L14_U1_xorInst_U4 ( .A(top_XOR_L14_U1_xorInst_n10), .ZN(
        top_XOR_L14_U1_xorInst_n11) );
  OR2_X1 top_XOR_L14_U1_xorInst_U3 ( .A1(top_XOR_L14_U1_xorInst_n9), .A2(
        Fresh[22]), .ZN(top_XOR_L14_U1_xorInst_n10) );
  AND2_X1 top_XOR_L14_U1_xorInst_U2 ( .A1(Fresh[22]), .A2(
        top_XOR_L14_U1_xorInst_n9), .ZN(top_XOR_L14_U1_xorInst_n12) );
  INV_X1 top_XOR_L14_U1_xorInst_U1 ( .A(Fresh[31]), .ZN(
        top_XOR_L14_U1_xorInst_n9) );
  AND2_X1 top_XOR_L14_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_343), .A2(
        top_new_AGEMA_signal_336), .ZN(top_XOR_L14_U1_w[0]) );
  AND2_X1 top_XOR_L14_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_344), .A2(
        top_new_AGEMA_signal_335), .ZN(top_XOR_L14_U1_w[1]) );
  AND2_X1 top_XOR_L14_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_344), .A2(
        top_new_AGEMA_signal_336), .ZN(top_XOR_L14_U1_w[2]) );
  AND2_X1 top_XOR_L14_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_343), .A2(
        top_new_AGEMA_signal_335), .ZN(top_XOR_L14_U1_w[3]) );
  OR2_X1 top_XOR_L14_U1_orInst1_U1 ( .A1(top_XOR_L14_U1_w[0]), .A2(
        top_XOR_L14_U1_w[1]), .ZN(top_new_AGEMA_signal_365) );
  OR2_X1 top_XOR_L14_U1_orInst2_U1 ( .A1(top_XOR_L14_U1_w[2]), .A2(
        top_XOR_L14_U1_w[3]), .ZN(top_new_AGEMA_signal_366) );
  OR2_X1 top_XOR_L15_U1_xorInst_U5 ( .A1(top_XOR_L15_U1_xorInst_n12), .A2(
        top_XOR_L15_U1_xorInst_n11), .ZN(top_L15) );
  INV_X1 top_XOR_L15_U1_xorInst_U4 ( .A(top_XOR_L15_U1_xorInst_n10), .ZN(
        top_XOR_L15_U1_xorInst_n11) );
  OR2_X1 top_XOR_L15_U1_xorInst_U3 ( .A1(top_XOR_L15_U1_xorInst_n9), .A2(
        Fresh[25]), .ZN(top_XOR_L15_U1_xorInst_n10) );
  AND2_X1 top_XOR_L15_U1_xorInst_U2 ( .A1(Fresh[25]), .A2(
        top_XOR_L15_U1_xorInst_n9), .ZN(top_XOR_L15_U1_xorInst_n12) );
  INV_X1 top_XOR_L15_U1_xorInst_U1 ( .A(top_L1), .ZN(top_XOR_L15_U1_xorInst_n9) );
  AND2_X1 top_XOR_L15_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_347), .A2(
        top_new_AGEMA_signal_340), .ZN(top_XOR_L15_U1_w[0]) );
  AND2_X1 top_XOR_L15_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_348), .A2(
        top_new_AGEMA_signal_339), .ZN(top_XOR_L15_U1_w[1]) );
  AND2_X1 top_XOR_L15_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_348), .A2(
        top_new_AGEMA_signal_340), .ZN(top_XOR_L15_U1_w[2]) );
  AND2_X1 top_XOR_L15_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_347), .A2(
        top_new_AGEMA_signal_339), .ZN(top_XOR_L15_U1_w[3]) );
  OR2_X1 top_XOR_L15_U1_orInst1_U1 ( .A1(top_XOR_L15_U1_w[0]), .A2(
        top_XOR_L15_U1_w[1]), .ZN(top_new_AGEMA_signal_367) );
  OR2_X1 top_XOR_L15_U1_orInst2_U1 ( .A1(top_XOR_L15_U1_w[2]), .A2(
        top_XOR_L15_U1_w[3]), .ZN(top_new_AGEMA_signal_368) );
  OR2_X1 top_XOR_L16_U1_xorInst_U5 ( .A1(top_XOR_L16_U1_xorInst_n12), .A2(
        top_XOR_L16_U1_xorInst_n11), .ZN(top_L16) );
  INV_X1 top_XOR_L16_U1_xorInst_U4 ( .A(top_XOR_L16_U1_xorInst_n10), .ZN(
        top_XOR_L16_U1_xorInst_n11) );
  OR2_X1 top_XOR_L16_U1_xorInst_U3 ( .A1(top_XOR_L16_U1_xorInst_n9), .A2(
        Fresh[26]), .ZN(top_XOR_L16_U1_xorInst_n10) );
  AND2_X1 top_XOR_L16_U1_xorInst_U2 ( .A1(Fresh[26]), .A2(
        top_XOR_L16_U1_xorInst_n9), .ZN(top_XOR_L16_U1_xorInst_n12) );
  INV_X1 top_XOR_L16_U1_xorInst_U1 ( .A(top_L0), .ZN(top_XOR_L16_U1_xorInst_n9) );
  AND2_X1 top_XOR_L16_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_373), .A2(
        top_new_AGEMA_signal_322), .ZN(top_XOR_L16_U1_w[0]) );
  AND2_X1 top_XOR_L16_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_374), .A2(
        top_new_AGEMA_signal_321), .ZN(top_XOR_L16_U1_w[1]) );
  AND2_X1 top_XOR_L16_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_374), .A2(
        top_new_AGEMA_signal_322), .ZN(top_XOR_L16_U1_w[2]) );
  AND2_X1 top_XOR_L16_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_373), .A2(
        top_new_AGEMA_signal_321), .ZN(top_XOR_L16_U1_w[3]) );
  OR2_X1 top_XOR_L16_U1_orInst1_U1 ( .A1(top_XOR_L16_U1_w[0]), .A2(
        top_XOR_L16_U1_w[1]), .ZN(top_new_AGEMA_signal_393) );
  OR2_X1 top_XOR_L16_U1_orInst2_U1 ( .A1(top_XOR_L16_U1_w[2]), .A2(
        top_XOR_L16_U1_w[3]), .ZN(top_new_AGEMA_signal_394) );
  OR2_X1 top_XOR_L17_U1_xorInst_U5 ( .A1(top_XOR_L17_U1_xorInst_n12), .A2(
        top_XOR_L17_U1_xorInst_n11), .ZN(top_L17) );
  INV_X1 top_XOR_L17_U1_xorInst_U4 ( .A(top_XOR_L17_U1_xorInst_n10), .ZN(
        top_XOR_L17_U1_xorInst_n11) );
  OR2_X1 top_XOR_L17_U1_xorInst_U3 ( .A1(top_XOR_L17_U1_xorInst_n9), .A2(
        Fresh[27]), .ZN(top_XOR_L17_U1_xorInst_n10) );
  AND2_X1 top_XOR_L17_U1_xorInst_U2 ( .A1(Fresh[27]), .A2(
        top_XOR_L17_U1_xorInst_n9), .ZN(top_XOR_L17_U1_xorInst_n12) );
  INV_X1 top_XOR_L17_U1_xorInst_U1 ( .A(top_L1), .ZN(top_XOR_L17_U1_xorInst_n9) );
  AND2_X1 top_XOR_L17_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_347), .A2(
        top_new_AGEMA_signal_324), .ZN(top_XOR_L17_U1_w[0]) );
  AND2_X1 top_XOR_L17_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_348), .A2(
        top_new_AGEMA_signal_323), .ZN(top_XOR_L17_U1_w[1]) );
  AND2_X1 top_XOR_L17_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_348), .A2(
        top_new_AGEMA_signal_324), .ZN(top_XOR_L17_U1_w[2]) );
  AND2_X1 top_XOR_L17_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_347), .A2(
        top_new_AGEMA_signal_323), .ZN(top_XOR_L17_U1_w[3]) );
  OR2_X1 top_XOR_L17_U1_orInst1_U1 ( .A1(top_XOR_L17_U1_w[0]), .A2(
        top_XOR_L17_U1_w[1]), .ZN(top_new_AGEMA_signal_369) );
  OR2_X1 top_XOR_L17_U1_orInst2_U1 ( .A1(top_XOR_L17_U1_w[2]), .A2(
        top_XOR_L17_U1_w[3]), .ZN(top_new_AGEMA_signal_370) );
  OR2_X1 top_XOR_L18_U1_xorInst_U5 ( .A1(top_XOR_L18_U1_xorInst_n12), .A2(
        top_XOR_L18_U1_xorInst_n11), .ZN(top_L18) );
  INV_X1 top_XOR_L18_U1_xorInst_U4 ( .A(top_XOR_L18_U1_xorInst_n10), .ZN(
        top_XOR_L18_U1_xorInst_n11) );
  OR2_X1 top_XOR_L18_U1_xorInst_U3 ( .A1(top_XOR_L18_U1_xorInst_n9), .A2(
        Fresh[28]), .ZN(top_XOR_L18_U1_xorInst_n10) );
  AND2_X1 top_XOR_L18_U1_xorInst_U2 ( .A1(Fresh[28]), .A2(
        top_XOR_L18_U1_xorInst_n9), .ZN(top_XOR_L18_U1_xorInst_n12) );
  INV_X1 top_XOR_L18_U1_xorInst_U1 ( .A(top_L8), .ZN(top_XOR_L18_U1_xorInst_n9) );
  AND2_X1 top_XOR_L18_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_349), .A2(
        top_new_AGEMA_signal_342), .ZN(top_XOR_L18_U1_w[0]) );
  AND2_X1 top_XOR_L18_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_350), .A2(
        top_new_AGEMA_signal_341), .ZN(top_XOR_L18_U1_w[1]) );
  AND2_X1 top_XOR_L18_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_350), .A2(
        top_new_AGEMA_signal_342), .ZN(top_XOR_L18_U1_w[2]) );
  AND2_X1 top_XOR_L18_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_349), .A2(
        top_new_AGEMA_signal_341), .ZN(top_XOR_L18_U1_w[3]) );
  OR2_X1 top_XOR_L18_U1_orInst1_U1 ( .A1(top_XOR_L18_U1_w[0]), .A2(
        top_XOR_L18_U1_w[1]), .ZN(top_new_AGEMA_signal_371) );
  OR2_X1 top_XOR_L18_U1_orInst2_U1 ( .A1(top_XOR_L18_U1_w[2]), .A2(
        top_XOR_L18_U1_w[3]), .ZN(top_new_AGEMA_signal_372) );
  OR2_X1 top_XOR_L19_U1_xorInst_U5 ( .A1(top_XOR_L19_U1_xorInst_n12), .A2(
        top_XOR_L19_U1_xorInst_n11), .ZN(top_L19) );
  INV_X1 top_XOR_L19_U1_xorInst_U4 ( .A(top_XOR_L19_U1_xorInst_n10), .ZN(
        top_XOR_L19_U1_xorInst_n11) );
  OR2_X1 top_XOR_L19_U1_xorInst_U3 ( .A1(top_XOR_L19_U1_xorInst_n9), .A2(
        Fresh[33]), .ZN(top_XOR_L19_U1_xorInst_n10) );
  AND2_X1 top_XOR_L19_U1_xorInst_U2 ( .A1(Fresh[33]), .A2(
        top_XOR_L19_U1_xorInst_n9), .ZN(top_XOR_L19_U1_xorInst_n12) );
  INV_X1 top_XOR_L19_U1_xorInst_U1 ( .A(top_L4), .ZN(top_XOR_L19_U1_xorInst_n9) );
  AND2_X1 top_XOR_L19_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_361), .A2(
        top_new_AGEMA_signal_346), .ZN(top_XOR_L19_U1_w[0]) );
  AND2_X1 top_XOR_L19_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_362), .A2(
        top_new_AGEMA_signal_345), .ZN(top_XOR_L19_U1_w[1]) );
  AND2_X1 top_XOR_L19_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_362), .A2(
        top_new_AGEMA_signal_346), .ZN(top_XOR_L19_U1_w[2]) );
  AND2_X1 top_XOR_L19_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_361), .A2(
        top_new_AGEMA_signal_345), .ZN(top_XOR_L19_U1_w[3]) );
  OR2_X1 top_XOR_L19_U1_orInst1_U1 ( .A1(top_XOR_L19_U1_w[0]), .A2(
        top_XOR_L19_U1_w[1]), .ZN(top_new_AGEMA_signal_385) );
  OR2_X1 top_XOR_L19_U1_orInst2_U1 ( .A1(top_XOR_L19_U1_w[2]), .A2(
        top_XOR_L19_U1_w[3]), .ZN(top_new_AGEMA_signal_386) );
  OR2_X1 top_XOR_L20_U1_xorInst_U5 ( .A1(top_XOR_L20_U1_xorInst_n12), .A2(
        top_XOR_L20_U1_xorInst_n11), .ZN(top_L20) );
  INV_X1 top_XOR_L20_U1_xorInst_U4 ( .A(top_XOR_L20_U1_xorInst_n10), .ZN(
        top_XOR_L20_U1_xorInst_n11) );
  OR2_X1 top_XOR_L20_U1_xorInst_U3 ( .A1(top_XOR_L20_U1_xorInst_n9), .A2(
        top_L0), .ZN(top_XOR_L20_U1_xorInst_n10) );
  AND2_X1 top_XOR_L20_U1_xorInst_U2 ( .A1(top_L0), .A2(
        top_XOR_L20_U1_xorInst_n9), .ZN(top_XOR_L20_U1_xorInst_n12) );
  INV_X1 top_XOR_L20_U1_xorInst_U1 ( .A(top_L1), .ZN(top_XOR_L20_U1_xorInst_n9) );
  AND2_X1 top_XOR_L20_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_347), .A2(
        top_new_AGEMA_signal_374), .ZN(top_XOR_L20_U1_w[0]) );
  AND2_X1 top_XOR_L20_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_348), .A2(
        top_new_AGEMA_signal_373), .ZN(top_XOR_L20_U1_w[1]) );
  AND2_X1 top_XOR_L20_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_348), .A2(
        top_new_AGEMA_signal_374), .ZN(top_XOR_L20_U1_w[2]) );
  AND2_X1 top_XOR_L20_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_347), .A2(
        top_new_AGEMA_signal_373), .ZN(top_XOR_L20_U1_w[3]) );
  OR2_X1 top_XOR_L20_U1_orInst1_U1 ( .A1(top_XOR_L20_U1_w[0]), .A2(
        top_XOR_L20_U1_w[1]), .ZN(top_new_AGEMA_signal_395) );
  OR2_X1 top_XOR_L20_U1_orInst2_U1 ( .A1(top_XOR_L20_U1_w[2]), .A2(
        top_XOR_L20_U1_w[3]), .ZN(top_new_AGEMA_signal_396) );
  OR2_X1 top_XOR_L21_U1_xorInst_U5 ( .A1(top_XOR_L21_U1_xorInst_n12), .A2(
        top_XOR_L21_U1_xorInst_n11), .ZN(top_L21) );
  INV_X1 top_XOR_L21_U1_xorInst_U4 ( .A(top_XOR_L21_U1_xorInst_n10), .ZN(
        top_XOR_L21_U1_xorInst_n11) );
  OR2_X1 top_XOR_L21_U1_xorInst_U3 ( .A1(top_XOR_L21_U1_xorInst_n9), .A2(
        top_L1), .ZN(top_XOR_L21_U1_xorInst_n10) );
  AND2_X1 top_XOR_L21_U1_xorInst_U2 ( .A1(top_L1), .A2(
        top_XOR_L21_U1_xorInst_n9), .ZN(top_XOR_L21_U1_xorInst_n12) );
  INV_X1 top_XOR_L21_U1_xorInst_U1 ( .A(top_L7), .ZN(top_XOR_L21_U1_xorInst_n9) );
  AND2_X1 top_XOR_L21_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_377), .A2(
        top_new_AGEMA_signal_348), .ZN(top_XOR_L21_U1_w[0]) );
  AND2_X1 top_XOR_L21_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_378), .A2(
        top_new_AGEMA_signal_347), .ZN(top_XOR_L21_U1_w[1]) );
  AND2_X1 top_XOR_L21_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_378), .A2(
        top_new_AGEMA_signal_348), .ZN(top_XOR_L21_U1_w[2]) );
  AND2_X1 top_XOR_L21_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_377), .A2(
        top_new_AGEMA_signal_347), .ZN(top_XOR_L21_U1_w[3]) );
  OR2_X1 top_XOR_L21_U1_orInst1_U1 ( .A1(top_XOR_L21_U1_w[0]), .A2(
        top_XOR_L21_U1_w[1]), .ZN(top_new_AGEMA_signal_397) );
  OR2_X1 top_XOR_L21_U1_orInst2_U1 ( .A1(top_XOR_L21_U1_w[2]), .A2(
        top_XOR_L21_U1_w[3]), .ZN(top_new_AGEMA_signal_398) );
  OR2_X1 top_XOR_L22_U1_xorInst_U5 ( .A1(top_XOR_L22_U1_xorInst_n12), .A2(
        top_XOR_L22_U1_xorInst_n11), .ZN(top_L22) );
  INV_X1 top_XOR_L22_U1_xorInst_U4 ( .A(top_XOR_L22_U1_xorInst_n10), .ZN(
        top_XOR_L22_U1_xorInst_n11) );
  OR2_X1 top_XOR_L22_U1_xorInst_U3 ( .A1(top_XOR_L22_U1_xorInst_n9), .A2(
        top_L3), .ZN(top_XOR_L22_U1_xorInst_n10) );
  AND2_X1 top_XOR_L22_U1_xorInst_U2 ( .A1(top_L3), .A2(
        top_XOR_L22_U1_xorInst_n9), .ZN(top_XOR_L22_U1_xorInst_n12) );
  INV_X1 top_XOR_L22_U1_xorInst_U1 ( .A(top_L12), .ZN(
        top_XOR_L22_U1_xorInst_n9) );
  AND2_X1 top_XOR_L22_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_351), .A2(
        top_new_AGEMA_signal_360), .ZN(top_XOR_L22_U1_w[0]) );
  AND2_X1 top_XOR_L22_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_352), .A2(
        top_new_AGEMA_signal_359), .ZN(top_XOR_L22_U1_w[1]) );
  AND2_X1 top_XOR_L22_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_352), .A2(
        top_new_AGEMA_signal_360), .ZN(top_XOR_L22_U1_w[2]) );
  AND2_X1 top_XOR_L22_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_351), .A2(
        top_new_AGEMA_signal_359), .ZN(top_XOR_L22_U1_w[3]) );
  OR2_X1 top_XOR_L22_U1_orInst1_U1 ( .A1(top_XOR_L22_U1_w[0]), .A2(
        top_XOR_L22_U1_w[1]), .ZN(top_new_AGEMA_signal_387) );
  OR2_X1 top_XOR_L22_U1_orInst2_U1 ( .A1(top_XOR_L22_U1_w[2]), .A2(
        top_XOR_L22_U1_w[3]), .ZN(top_new_AGEMA_signal_388) );
  OR2_X1 top_XOR_L23_U1_xorInst_U5 ( .A1(top_XOR_L23_U1_xorInst_n12), .A2(
        top_XOR_L23_U1_xorInst_n11), .ZN(top_L23) );
  INV_X1 top_XOR_L23_U1_xorInst_U4 ( .A(top_XOR_L23_U1_xorInst_n10), .ZN(
        top_XOR_L23_U1_xorInst_n11) );
  OR2_X1 top_XOR_L23_U1_xorInst_U3 ( .A1(top_XOR_L23_U1_xorInst_n9), .A2(
        top_L18), .ZN(top_XOR_L23_U1_xorInst_n10) );
  AND2_X1 top_XOR_L23_U1_xorInst_U2 ( .A1(top_L18), .A2(
        top_XOR_L23_U1_xorInst_n9), .ZN(top_XOR_L23_U1_xorInst_n12) );
  INV_X1 top_XOR_L23_U1_xorInst_U1 ( .A(top_L2), .ZN(top_XOR_L23_U1_xorInst_n9) );
  AND2_X1 top_XOR_L23_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_357), .A2(
        top_new_AGEMA_signal_372), .ZN(top_XOR_L23_U1_w[0]) );
  AND2_X1 top_XOR_L23_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_358), .A2(
        top_new_AGEMA_signal_371), .ZN(top_XOR_L23_U1_w[1]) );
  AND2_X1 top_XOR_L23_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_358), .A2(
        top_new_AGEMA_signal_372), .ZN(top_XOR_L23_U1_w[2]) );
  AND2_X1 top_XOR_L23_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_357), .A2(
        top_new_AGEMA_signal_371), .ZN(top_XOR_L23_U1_w[3]) );
  OR2_X1 top_XOR_L23_U1_orInst1_U1 ( .A1(top_XOR_L23_U1_w[0]), .A2(
        top_XOR_L23_U1_w[1]), .ZN(top_new_AGEMA_signal_389) );
  OR2_X1 top_XOR_L23_U1_orInst2_U1 ( .A1(top_XOR_L23_U1_w[2]), .A2(
        top_XOR_L23_U1_w[3]), .ZN(top_new_AGEMA_signal_390) );
  OR2_X1 top_XOR_L24_U1_xorInst_U5 ( .A1(top_XOR_L24_U1_xorInst_n12), .A2(
        top_XOR_L24_U1_xorInst_n11), .ZN(top_L24) );
  INV_X1 top_XOR_L24_U1_xorInst_U4 ( .A(top_XOR_L24_U1_xorInst_n10), .ZN(
        top_XOR_L24_U1_xorInst_n11) );
  OR2_X1 top_XOR_L24_U1_xorInst_U3 ( .A1(top_XOR_L24_U1_xorInst_n9), .A2(
        top_L15), .ZN(top_XOR_L24_U1_xorInst_n10) );
  AND2_X1 top_XOR_L24_U1_xorInst_U2 ( .A1(top_L15), .A2(
        top_XOR_L24_U1_xorInst_n9), .ZN(top_XOR_L24_U1_xorInst_n12) );
  INV_X1 top_XOR_L24_U1_xorInst_U1 ( .A(top_L9), .ZN(top_XOR_L24_U1_xorInst_n9) );
  AND2_X1 top_XOR_L24_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_379), .A2(
        top_new_AGEMA_signal_368), .ZN(top_XOR_L24_U1_w[0]) );
  AND2_X1 top_XOR_L24_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_380), .A2(
        top_new_AGEMA_signal_367), .ZN(top_XOR_L24_U1_w[1]) );
  AND2_X1 top_XOR_L24_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_380), .A2(
        top_new_AGEMA_signal_368), .ZN(top_XOR_L24_U1_w[2]) );
  AND2_X1 top_XOR_L24_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_379), .A2(
        top_new_AGEMA_signal_367), .ZN(top_XOR_L24_U1_w[3]) );
  OR2_X1 top_XOR_L24_U1_orInst1_U1 ( .A1(top_XOR_L24_U1_w[0]), .A2(
        top_XOR_L24_U1_w[1]), .ZN(top_new_AGEMA_signal_399) );
  OR2_X1 top_XOR_L24_U1_orInst2_U1 ( .A1(top_XOR_L24_U1_w[2]), .A2(
        top_XOR_L24_U1_w[3]), .ZN(top_new_AGEMA_signal_400) );
  OR2_X1 top_XOR_L25_U1_xorInst_U5 ( .A1(top_XOR_L25_U1_xorInst_n12), .A2(
        top_XOR_L25_U1_xorInst_n11), .ZN(top_L25) );
  INV_X1 top_XOR_L25_U1_xorInst_U4 ( .A(top_XOR_L25_U1_xorInst_n10), .ZN(
        top_XOR_L25_U1_xorInst_n11) );
  OR2_X1 top_XOR_L25_U1_xorInst_U3 ( .A1(top_XOR_L25_U1_xorInst_n9), .A2(
        top_L6), .ZN(top_XOR_L25_U1_xorInst_n10) );
  AND2_X1 top_XOR_L25_U1_xorInst_U2 ( .A1(top_L6), .A2(
        top_XOR_L25_U1_xorInst_n9), .ZN(top_XOR_L25_U1_xorInst_n12) );
  INV_X1 top_XOR_L25_U1_xorInst_U1 ( .A(top_L10), .ZN(
        top_XOR_L25_U1_xorInst_n9) );
  AND2_X1 top_XOR_L25_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_381), .A2(
        top_new_AGEMA_signal_376), .ZN(top_XOR_L25_U1_w[0]) );
  AND2_X1 top_XOR_L25_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_382), .A2(
        top_new_AGEMA_signal_375), .ZN(top_XOR_L25_U1_w[1]) );
  AND2_X1 top_XOR_L25_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_382), .A2(
        top_new_AGEMA_signal_376), .ZN(top_XOR_L25_U1_w[2]) );
  AND2_X1 top_XOR_L25_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_381), .A2(
        top_new_AGEMA_signal_375), .ZN(top_XOR_L25_U1_w[3]) );
  OR2_X1 top_XOR_L25_U1_orInst1_U1 ( .A1(top_XOR_L25_U1_w[0]), .A2(
        top_XOR_L25_U1_w[1]), .ZN(top_new_AGEMA_signal_401) );
  OR2_X1 top_XOR_L25_U1_orInst2_U1 ( .A1(top_XOR_L25_U1_w[2]), .A2(
        top_XOR_L25_U1_w[3]), .ZN(top_new_AGEMA_signal_402) );
  OR2_X1 top_XOR_L26_U1_xorInst_U5 ( .A1(top_XOR_L26_U1_xorInst_n12), .A2(
        top_XOR_L26_U1_xorInst_n11), .ZN(top_L26) );
  INV_X1 top_XOR_L26_U1_xorInst_U4 ( .A(top_XOR_L26_U1_xorInst_n10), .ZN(
        top_XOR_L26_U1_xorInst_n11) );
  OR2_X1 top_XOR_L26_U1_xorInst_U3 ( .A1(top_XOR_L26_U1_xorInst_n9), .A2(
        top_L7), .ZN(top_XOR_L26_U1_xorInst_n10) );
  AND2_X1 top_XOR_L26_U1_xorInst_U2 ( .A1(top_L7), .A2(
        top_XOR_L26_U1_xorInst_n9), .ZN(top_XOR_L26_U1_xorInst_n12) );
  INV_X1 top_XOR_L26_U1_xorInst_U1 ( .A(top_L9), .ZN(top_XOR_L26_U1_xorInst_n9) );
  AND2_X1 top_XOR_L26_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_379), .A2(
        top_new_AGEMA_signal_378), .ZN(top_XOR_L26_U1_w[0]) );
  AND2_X1 top_XOR_L26_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_380), .A2(
        top_new_AGEMA_signal_377), .ZN(top_XOR_L26_U1_w[1]) );
  AND2_X1 top_XOR_L26_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_380), .A2(
        top_new_AGEMA_signal_378), .ZN(top_XOR_L26_U1_w[2]) );
  AND2_X1 top_XOR_L26_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_379), .A2(
        top_new_AGEMA_signal_377), .ZN(top_XOR_L26_U1_w[3]) );
  OR2_X1 top_XOR_L26_U1_orInst1_U1 ( .A1(top_XOR_L26_U1_w[0]), .A2(
        top_XOR_L26_U1_w[1]), .ZN(top_new_AGEMA_signal_403) );
  OR2_X1 top_XOR_L26_U1_orInst2_U1 ( .A1(top_XOR_L26_U1_w[2]), .A2(
        top_XOR_L26_U1_w[3]), .ZN(top_new_AGEMA_signal_404) );
  OR2_X1 top_XOR_L27_U1_xorInst_U5 ( .A1(top_XOR_L27_U1_xorInst_n12), .A2(
        top_XOR_L27_U1_xorInst_n11), .ZN(top_L27) );
  INV_X1 top_XOR_L27_U1_xorInst_U4 ( .A(top_XOR_L27_U1_xorInst_n10), .ZN(
        top_XOR_L27_U1_xorInst_n11) );
  OR2_X1 top_XOR_L27_U1_xorInst_U3 ( .A1(top_XOR_L27_U1_xorInst_n9), .A2(
        top_L8), .ZN(top_XOR_L27_U1_xorInst_n10) );
  AND2_X1 top_XOR_L27_U1_xorInst_U2 ( .A1(top_L8), .A2(
        top_XOR_L27_U1_xorInst_n9), .ZN(top_XOR_L27_U1_xorInst_n12) );
  INV_X1 top_XOR_L27_U1_xorInst_U1 ( .A(top_L10), .ZN(
        top_XOR_L27_U1_xorInst_n9) );
  AND2_X1 top_XOR_L27_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_381), .A2(
        top_new_AGEMA_signal_350), .ZN(top_XOR_L27_U1_w[0]) );
  AND2_X1 top_XOR_L27_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_382), .A2(
        top_new_AGEMA_signal_349), .ZN(top_XOR_L27_U1_w[1]) );
  AND2_X1 top_XOR_L27_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_382), .A2(
        top_new_AGEMA_signal_350), .ZN(top_XOR_L27_U1_w[2]) );
  AND2_X1 top_XOR_L27_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_381), .A2(
        top_new_AGEMA_signal_349), .ZN(top_XOR_L27_U1_w[3]) );
  OR2_X1 top_XOR_L27_U1_orInst1_U1 ( .A1(top_XOR_L27_U1_w[0]), .A2(
        top_XOR_L27_U1_w[1]), .ZN(top_new_AGEMA_signal_405) );
  OR2_X1 top_XOR_L27_U1_orInst2_U1 ( .A1(top_XOR_L27_U1_w[2]), .A2(
        top_XOR_L27_U1_w[3]), .ZN(top_new_AGEMA_signal_406) );
  OR2_X1 top_XOR_L28_U1_xorInst_U5 ( .A1(top_XOR_L28_U1_xorInst_n12), .A2(
        top_XOR_L28_U1_xorInst_n11), .ZN(top_L28) );
  INV_X1 top_XOR_L28_U1_xorInst_U4 ( .A(top_XOR_L28_U1_xorInst_n10), .ZN(
        top_XOR_L28_U1_xorInst_n11) );
  OR2_X1 top_XOR_L28_U1_xorInst_U3 ( .A1(top_XOR_L28_U1_xorInst_n9), .A2(
        top_L11), .ZN(top_XOR_L28_U1_xorInst_n10) );
  AND2_X1 top_XOR_L28_U1_xorInst_U2 ( .A1(top_L11), .A2(
        top_XOR_L28_U1_xorInst_n9), .ZN(top_XOR_L28_U1_xorInst_n12) );
  INV_X1 top_XOR_L28_U1_xorInst_U1 ( .A(top_L14), .ZN(
        top_XOR_L28_U1_xorInst_n9) );
  AND2_X1 top_XOR_L28_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_365), .A2(
        top_new_AGEMA_signal_384), .ZN(top_XOR_L28_U1_w[0]) );
  AND2_X1 top_XOR_L28_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_366), .A2(
        top_new_AGEMA_signal_383), .ZN(top_XOR_L28_U1_w[1]) );
  AND2_X1 top_XOR_L28_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_366), .A2(
        top_new_AGEMA_signal_384), .ZN(top_XOR_L28_U1_w[2]) );
  AND2_X1 top_XOR_L28_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_365), .A2(
        top_new_AGEMA_signal_383), .ZN(top_XOR_L28_U1_w[3]) );
  OR2_X1 top_XOR_L28_U1_orInst1_U1 ( .A1(top_XOR_L28_U1_w[0]), .A2(
        top_XOR_L28_U1_w[1]), .ZN(top_new_AGEMA_signal_407) );
  OR2_X1 top_XOR_L28_U1_orInst2_U1 ( .A1(top_XOR_L28_U1_w[2]), .A2(
        top_XOR_L28_U1_w[3]), .ZN(top_new_AGEMA_signal_408) );
  OR2_X1 top_XOR_L29_U1_xorInst_U5 ( .A1(top_XOR_L29_U1_xorInst_n12), .A2(
        top_XOR_L29_U1_xorInst_n11), .ZN(top_L29) );
  INV_X1 top_XOR_L29_U1_xorInst_U4 ( .A(top_XOR_L29_U1_xorInst_n10), .ZN(
        top_XOR_L29_U1_xorInst_n11) );
  OR2_X1 top_XOR_L29_U1_xorInst_U3 ( .A1(top_XOR_L29_U1_xorInst_n9), .A2(
        top_L11), .ZN(top_XOR_L29_U1_xorInst_n10) );
  AND2_X1 top_XOR_L29_U1_xorInst_U2 ( .A1(top_L11), .A2(
        top_XOR_L29_U1_xorInst_n9), .ZN(top_XOR_L29_U1_xorInst_n12) );
  INV_X1 top_XOR_L29_U1_xorInst_U1 ( .A(top_L17), .ZN(
        top_XOR_L29_U1_xorInst_n9) );
  AND2_X1 top_XOR_L29_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_369), .A2(
        top_new_AGEMA_signal_384), .ZN(top_XOR_L29_U1_w[0]) );
  AND2_X1 top_XOR_L29_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_370), .A2(
        top_new_AGEMA_signal_383), .ZN(top_XOR_L29_U1_w[1]) );
  AND2_X1 top_XOR_L29_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_370), .A2(
        top_new_AGEMA_signal_384), .ZN(top_XOR_L29_U1_w[2]) );
  AND2_X1 top_XOR_L29_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_369), .A2(
        top_new_AGEMA_signal_383), .ZN(top_XOR_L29_U1_w[3]) );
  OR2_X1 top_XOR_L29_U1_orInst1_U1 ( .A1(top_XOR_L29_U1_w[0]), .A2(
        top_XOR_L29_U1_w[1]), .ZN(top_new_AGEMA_signal_409) );
  OR2_X1 top_XOR_L29_U1_orInst2_U1 ( .A1(top_XOR_L29_U1_w[2]), .A2(
        top_XOR_L29_U1_w[3]), .ZN(top_new_AGEMA_signal_410) );
  OR2_X1 top_XOR_S0_U1_xorInst_U5 ( .A1(top_XOR_S0_U1_xorInst_n12), .A2(
        top_XOR_S0_U1_xorInst_n11), .ZN(Y_s0[7]) );
  INV_X1 top_XOR_S0_U1_xorInst_U4 ( .A(top_XOR_S0_U1_xorInst_n10), .ZN(
        top_XOR_S0_U1_xorInst_n11) );
  OR2_X1 top_XOR_S0_U1_xorInst_U3 ( .A1(top_XOR_S0_U1_xorInst_n9), .A2(top_L6), 
        .ZN(top_XOR_S0_U1_xorInst_n10) );
  AND2_X1 top_XOR_S0_U1_xorInst_U2 ( .A1(top_L6), .A2(top_XOR_S0_U1_xorInst_n9), .ZN(top_XOR_S0_U1_xorInst_n12) );
  INV_X1 top_XOR_S0_U1_xorInst_U1 ( .A(top_L24), .ZN(top_XOR_S0_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_S0_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_399), .A2(
        top_new_AGEMA_signal_376), .ZN(top_XOR_S0_U1_w[0]) );
  AND2_X1 top_XOR_S0_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_400), .A2(
        top_new_AGEMA_signal_375), .ZN(top_XOR_S0_U1_w[1]) );
  AND2_X1 top_XOR_S0_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_400), .A2(
        top_new_AGEMA_signal_376), .ZN(top_XOR_S0_U1_w[2]) );
  AND2_X1 top_XOR_S0_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_399), .A2(
        top_new_AGEMA_signal_375), .ZN(top_XOR_S0_U1_w[3]) );
  OR2_X1 top_XOR_S0_U1_orInst1_U1 ( .A1(top_XOR_S0_U1_w[0]), .A2(
        top_XOR_S0_U1_w[1]), .ZN(Y_s1[7]) );
  OR2_X1 top_XOR_S0_U1_orInst2_U1 ( .A1(top_XOR_S0_U1_w[2]), .A2(
        top_XOR_S0_U1_w[3]), .ZN(top_XOR_S0_U1_c_2_) );
  OR2_X1 top_XOR_S1_U1_xorInst_U5 ( .A1(top_XOR_S1_U1_xorInst_n12), .A2(
        top_XOR_S1_U1_xorInst_n11), .ZN(Y_s0[6]) );
  INV_X1 top_XOR_S1_U1_xorInst_U4 ( .A(top_XOR_S1_U1_xorInst_n10), .ZN(
        top_XOR_S1_U1_xorInst_n11) );
  OR2_X1 top_XOR_S1_U1_xorInst_U3 ( .A1(top_XOR_S1_U1_xorInst_n9), .A2(top_L16), .ZN(top_XOR_S1_U1_xorInst_n10) );
  AND2_X1 top_XOR_S1_U1_xorInst_U2 ( .A1(top_L16), .A2(
        top_XOR_S1_U1_xorInst_n9), .ZN(top_XOR_S1_U1_xorInst_n12) );
  INV_X1 top_XOR_S1_U1_xorInst_U1 ( .A(top_L26), .ZN(top_XOR_S1_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_S1_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_403), .A2(
        top_new_AGEMA_signal_394), .ZN(top_XOR_S1_U1_w[0]) );
  AND2_X1 top_XOR_S1_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_404), .A2(
        top_new_AGEMA_signal_393), .ZN(top_XOR_S1_U1_w[1]) );
  AND2_X1 top_XOR_S1_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_404), .A2(
        top_new_AGEMA_signal_394), .ZN(top_XOR_S1_U1_w[2]) );
  AND2_X1 top_XOR_S1_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_403), .A2(
        top_new_AGEMA_signal_393), .ZN(top_XOR_S1_U1_w[3]) );
  OR2_X1 top_XOR_S1_U1_orInst1_U1 ( .A1(top_XOR_S1_U1_w[0]), .A2(
        top_XOR_S1_U1_w[1]), .ZN(top_XOR_S1_U1_c_2_) );
  OR2_X1 top_XOR_S1_U1_orInst2_U1 ( .A1(top_XOR_S1_U1_w[2]), .A2(
        top_XOR_S1_U1_w[3]), .ZN(Y_s1[6]) );
  OR2_X1 top_XOR_S2_U1_xorInst_U5 ( .A1(top_XOR_S2_U1_xorInst_n12), .A2(
        top_XOR_S2_U1_xorInst_n11), .ZN(Y_s0[5]) );
  INV_X1 top_XOR_S2_U1_xorInst_U4 ( .A(top_XOR_S2_U1_xorInst_n10), .ZN(
        top_XOR_S2_U1_xorInst_n11) );
  OR2_X1 top_XOR_S2_U1_xorInst_U3 ( .A1(top_XOR_S2_U1_xorInst_n9), .A2(top_L19), .ZN(top_XOR_S2_U1_xorInst_n10) );
  AND2_X1 top_XOR_S2_U1_xorInst_U2 ( .A1(top_L19), .A2(
        top_XOR_S2_U1_xorInst_n9), .ZN(top_XOR_S2_U1_xorInst_n12) );
  INV_X1 top_XOR_S2_U1_xorInst_U1 ( .A(top_L28), .ZN(top_XOR_S2_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_S2_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_407), .A2(
        top_new_AGEMA_signal_386), .ZN(top_XOR_S2_U1_w[0]) );
  AND2_X1 top_XOR_S2_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_408), .A2(
        top_new_AGEMA_signal_385), .ZN(top_XOR_S2_U1_w[1]) );
  AND2_X1 top_XOR_S2_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_408), .A2(
        top_new_AGEMA_signal_386), .ZN(top_XOR_S2_U1_w[2]) );
  AND2_X1 top_XOR_S2_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_407), .A2(
        top_new_AGEMA_signal_385), .ZN(top_XOR_S2_U1_w[3]) );
  OR2_X1 top_XOR_S2_U1_orInst1_U1 ( .A1(top_XOR_S2_U1_w[0]), .A2(
        top_XOR_S2_U1_w[1]), .ZN(top_XOR_S2_U1_c_2_) );
  OR2_X1 top_XOR_S2_U1_orInst2_U1 ( .A1(top_XOR_S2_U1_w[2]), .A2(
        top_XOR_S2_U1_w[3]), .ZN(Y_s1[5]) );
  OR2_X1 top_XOR_S3_U1_xorInst_U5 ( .A1(top_XOR_S3_U1_xorInst_n12), .A2(
        top_XOR_S3_U1_xorInst_n11), .ZN(Y_s0[4]) );
  INV_X1 top_XOR_S3_U1_xorInst_U4 ( .A(top_XOR_S3_U1_xorInst_n10), .ZN(
        top_XOR_S3_U1_xorInst_n11) );
  OR2_X1 top_XOR_S3_U1_xorInst_U3 ( .A1(top_XOR_S3_U1_xorInst_n9), .A2(top_L6), 
        .ZN(top_XOR_S3_U1_xorInst_n10) );
  AND2_X1 top_XOR_S3_U1_xorInst_U2 ( .A1(top_L6), .A2(top_XOR_S3_U1_xorInst_n9), .ZN(top_XOR_S3_U1_xorInst_n12) );
  INV_X1 top_XOR_S3_U1_xorInst_U1 ( .A(top_L21), .ZN(top_XOR_S3_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_S3_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_397), .A2(
        top_new_AGEMA_signal_376), .ZN(top_XOR_S3_U1_w[0]) );
  AND2_X1 top_XOR_S3_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_398), .A2(
        top_new_AGEMA_signal_375), .ZN(top_XOR_S3_U1_w[1]) );
  AND2_X1 top_XOR_S3_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_398), .A2(
        top_new_AGEMA_signal_376), .ZN(top_XOR_S3_U1_w[2]) );
  AND2_X1 top_XOR_S3_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_397), .A2(
        top_new_AGEMA_signal_375), .ZN(top_XOR_S3_U1_w[3]) );
  OR2_X1 top_XOR_S3_U1_orInst1_U1 ( .A1(top_XOR_S3_U1_w[0]), .A2(
        top_XOR_S3_U1_w[1]), .ZN(Y_s1[4]) );
  OR2_X1 top_XOR_S3_U1_orInst2_U1 ( .A1(top_XOR_S3_U1_w[2]), .A2(
        top_XOR_S3_U1_w[3]), .ZN(top_XOR_S3_U1_c_2_) );
  OR2_X1 top_XOR_S4_U1_xorInst_U5 ( .A1(top_XOR_S4_U1_xorInst_n12), .A2(
        top_XOR_S4_U1_xorInst_n11), .ZN(Y_s0[3]) );
  INV_X1 top_XOR_S4_U1_xorInst_U4 ( .A(top_XOR_S4_U1_xorInst_n10), .ZN(
        top_XOR_S4_U1_xorInst_n11) );
  OR2_X1 top_XOR_S4_U1_xorInst_U3 ( .A1(top_XOR_S4_U1_xorInst_n9), .A2(top_L20), .ZN(top_XOR_S4_U1_xorInst_n10) );
  AND2_X1 top_XOR_S4_U1_xorInst_U2 ( .A1(top_L20), .A2(
        top_XOR_S4_U1_xorInst_n9), .ZN(top_XOR_S4_U1_xorInst_n12) );
  INV_X1 top_XOR_S4_U1_xorInst_U1 ( .A(top_L22), .ZN(top_XOR_S4_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_S4_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_387), .A2(
        top_new_AGEMA_signal_396), .ZN(top_XOR_S4_U1_w[0]) );
  AND2_X1 top_XOR_S4_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_388), .A2(
        top_new_AGEMA_signal_395), .ZN(top_XOR_S4_U1_w[1]) );
  AND2_X1 top_XOR_S4_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_388), .A2(
        top_new_AGEMA_signal_396), .ZN(top_XOR_S4_U1_w[2]) );
  AND2_X1 top_XOR_S4_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_387), .A2(
        top_new_AGEMA_signal_395), .ZN(top_XOR_S4_U1_w[3]) );
  OR2_X1 top_XOR_S4_U1_orInst1_U1 ( .A1(top_XOR_S4_U1_w[0]), .A2(
        top_XOR_S4_U1_w[1]), .ZN(Y_s1[3]) );
  OR2_X1 top_XOR_S4_U1_orInst2_U1 ( .A1(top_XOR_S4_U1_w[2]), .A2(
        top_XOR_S4_U1_w[3]), .ZN(top_XOR_S4_U1_c_2_) );
  OR2_X1 top_XOR_S5_U1_xorInst_U5 ( .A1(top_XOR_S5_U1_xorInst_n12), .A2(
        top_XOR_S5_U1_xorInst_n11), .ZN(Y_s0[2]) );
  INV_X1 top_XOR_S5_U1_xorInst_U4 ( .A(top_XOR_S5_U1_xorInst_n10), .ZN(
        top_XOR_S5_U1_xorInst_n11) );
  OR2_X1 top_XOR_S5_U1_xorInst_U3 ( .A1(top_XOR_S5_U1_xorInst_n9), .A2(top_L25), .ZN(top_XOR_S5_U1_xorInst_n10) );
  AND2_X1 top_XOR_S5_U1_xorInst_U2 ( .A1(top_L25), .A2(
        top_XOR_S5_U1_xorInst_n9), .ZN(top_XOR_S5_U1_xorInst_n12) );
  INV_X1 top_XOR_S5_U1_xorInst_U1 ( .A(top_L29), .ZN(top_XOR_S5_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_S5_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_409), .A2(
        top_new_AGEMA_signal_402), .ZN(top_XOR_S5_U1_w[0]) );
  AND2_X1 top_XOR_S5_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_410), .A2(
        top_new_AGEMA_signal_401), .ZN(top_XOR_S5_U1_w[1]) );
  AND2_X1 top_XOR_S5_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_410), .A2(
        top_new_AGEMA_signal_402), .ZN(top_XOR_S5_U1_w[2]) );
  AND2_X1 top_XOR_S5_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_409), .A2(
        top_new_AGEMA_signal_401), .ZN(top_XOR_S5_U1_w[3]) );
  OR2_X1 top_XOR_S5_U1_orInst1_U1 ( .A1(top_XOR_S5_U1_w[0]), .A2(
        top_XOR_S5_U1_w[1]), .ZN(Y_s1[2]) );
  OR2_X1 top_XOR_S5_U1_orInst2_U1 ( .A1(top_XOR_S5_U1_w[2]), .A2(
        top_XOR_S5_U1_w[3]), .ZN(top_XOR_S5_U1_c_2_) );
  OR2_X1 top_XOR_S6_U1_xorInst_U5 ( .A1(top_XOR_S6_U1_xorInst_n12), .A2(
        top_XOR_S6_U1_xorInst_n11), .ZN(Y_s0[1]) );
  INV_X1 top_XOR_S6_U1_xorInst_U4 ( .A(top_XOR_S6_U1_xorInst_n10), .ZN(
        top_XOR_S6_U1_xorInst_n11) );
  OR2_X1 top_XOR_S6_U1_xorInst_U3 ( .A1(top_XOR_S6_U1_xorInst_n9), .A2(top_L13), .ZN(top_XOR_S6_U1_xorInst_n10) );
  AND2_X1 top_XOR_S6_U1_xorInst_U2 ( .A1(top_L13), .A2(
        top_XOR_S6_U1_xorInst_n9), .ZN(top_XOR_S6_U1_xorInst_n12) );
  INV_X1 top_XOR_S6_U1_xorInst_U1 ( .A(top_L27), .ZN(top_XOR_S6_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_S6_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_405), .A2(
        top_new_AGEMA_signal_392), .ZN(top_XOR_S6_U1_w[0]) );
  AND2_X1 top_XOR_S6_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_406), .A2(
        top_new_AGEMA_signal_391), .ZN(top_XOR_S6_U1_w[1]) );
  AND2_X1 top_XOR_S6_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_406), .A2(
        top_new_AGEMA_signal_392), .ZN(top_XOR_S6_U1_w[2]) );
  AND2_X1 top_XOR_S6_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_405), .A2(
        top_new_AGEMA_signal_391), .ZN(top_XOR_S6_U1_w[3]) );
  OR2_X1 top_XOR_S6_U1_orInst1_U1 ( .A1(top_XOR_S6_U1_w[0]), .A2(
        top_XOR_S6_U1_w[1]), .ZN(top_XOR_S6_U1_c_2_) );
  OR2_X1 top_XOR_S6_U1_orInst2_U1 ( .A1(top_XOR_S6_U1_w[2]), .A2(
        top_XOR_S6_U1_w[3]), .ZN(Y_s1[1]) );
  OR2_X1 top_XOR_S7_U1_xorInst_U5 ( .A1(top_XOR_S7_U1_xorInst_n12), .A2(
        top_XOR_S7_U1_xorInst_n11), .ZN(Y_s0[0]) );
  INV_X1 top_XOR_S7_U1_xorInst_U4 ( .A(top_XOR_S7_U1_xorInst_n10), .ZN(
        top_XOR_S7_U1_xorInst_n11) );
  OR2_X1 top_XOR_S7_U1_xorInst_U3 ( .A1(top_XOR_S7_U1_xorInst_n9), .A2(top_L6), 
        .ZN(top_XOR_S7_U1_xorInst_n10) );
  AND2_X1 top_XOR_S7_U1_xorInst_U2 ( .A1(top_L6), .A2(top_XOR_S7_U1_xorInst_n9), .ZN(top_XOR_S7_U1_xorInst_n12) );
  INV_X1 top_XOR_S7_U1_xorInst_U1 ( .A(top_L23), .ZN(top_XOR_S7_U1_xorInst_n9)
         );
  AND2_X1 top_XOR_S7_U1_andInst0_U1 ( .A1(top_new_AGEMA_signal_389), .A2(
        top_new_AGEMA_signal_376), .ZN(top_XOR_S7_U1_w[0]) );
  AND2_X1 top_XOR_S7_U1_andInst1_U1 ( .A1(top_new_AGEMA_signal_390), .A2(
        top_new_AGEMA_signal_375), .ZN(top_XOR_S7_U1_w[1]) );
  AND2_X1 top_XOR_S7_U1_andInst2_U1 ( .A1(top_new_AGEMA_signal_390), .A2(
        top_new_AGEMA_signal_376), .ZN(top_XOR_S7_U1_w[2]) );
  AND2_X1 top_XOR_S7_U1_andInst3_U1 ( .A1(top_new_AGEMA_signal_389), .A2(
        top_new_AGEMA_signal_375), .ZN(top_XOR_S7_U1_w[3]) );
  OR2_X1 top_XOR_S7_U1_orInst1_U1 ( .A1(top_XOR_S7_U1_w[0]), .A2(
        top_XOR_S7_U1_w[1]), .ZN(top_XOR_S7_U1_c_2_) );
  OR2_X1 top_XOR_S7_U1_orInst2_U1 ( .A1(top_XOR_S7_U1_w[2]), .A2(
        top_XOR_S7_U1_w[3]), .ZN(Y_s1[0]) );
endmodule

