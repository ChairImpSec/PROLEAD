module circuit ( ClkxCI, XxDI, Zmul1xDI, Zmul2xDI, Zmul3xDI, Zinv1xDI, 
        Zinv2xDI, Zinv3xDI, QxDO );
  input [31:0] XxDI;
  input [23:0] Zmul1xDI;
  input [23:0] Zmul2xDI;
  input [23:0] Zmul3xDI;
  input [11:0] Zinv1xDI;
  input [11:0] Zinv2xDI;
  input [11:0] Zinv3xDI;
  output [31:0] QxDO;
  input ClkxCI;
  wire   mappedxD_3__7_, mappedxD_3__6_, mappedxD_3__5_, mappedxD_3__4_,
         mappedxD_3__3_, mappedxD_3__1_, mappedxD_3__0_, mappedxD_2__7_,
         mappedxD_2__6_, mappedxD_2__5_, mappedxD_2__4_, mappedxD_2__3_,
         mappedxD_2__1_, mappedxD_2__0_, mappedxD_1__7_, mappedxD_1__6_,
         mappedxD_1__5_, mappedxD_1__4_, mappedxD_1__3_, mappedxD_1__1_,
         mappedxD_1__0_, mappedxD_0__7_, mappedxD_0__6_, mappedxD_0__5_,
         mappedxD_0__4_, mappedxD_0__3_, mappedxD_0__1_, mappedxD_0__0_,
         InvMappedxD_0__6_, InvMappedxD_0__5_, InvMappedxD_0__1_,
         InvMappedxD_0__0_, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, input_mapping_3_n23, input_mapping_3_n22,
         input_mapping_3_n21, input_mapping_3_n20, input_mapping_3_n19,
         input_mapping_3_n18, input_mapping_3_n17, output_mapping_3_n9,
         output_mapping_3_n8, output_mapping_3_n7, input_mapping_2_n23,
         input_mapping_2_n22, input_mapping_2_n21, input_mapping_2_n20,
         input_mapping_2_n19, input_mapping_2_n18, input_mapping_2_n17,
         output_mapping_2_n9, output_mapping_2_n8, output_mapping_2_n7,
         input_mapping_1_n23, input_mapping_1_n22, input_mapping_1_n21,
         input_mapping_1_n20, input_mapping_1_n19, input_mapping_1_n18,
         input_mapping_1_n17, output_mapping_1_n9, output_mapping_1_n8,
         output_mapping_1_n7, input_mapping_0_n23, input_mapping_0_n22,
         input_mapping_0_n21, input_mapping_0_n20, input_mapping_0_n19,
         input_mapping_0_n18, input_mapping_0_n17, output_mapping_0_n9,
         output_mapping_0_n8, output_mapping_0_n7, mul_y0y1_n32, mul_y0y1_n31,
         mul_y0y1_n30, mul_y0y1_n29, mul_y0y1_n28, mul_y0y1_n27, mul_y0y1_n26,
         mul_y0y1_n25, mul_y0y1_n24, mul_y0y1_n23, mul_y0y1_n22, mul_y0y1_n21,
         mul_y0y1_n20, mul_y0y1_n19, mul_y0y1_n18, mul_y0y1_n17, mul_y0y1_n16,
         mul_y0y1_n15, mul_y0y1_n14, mul_y0y1_n13, mul_y0y1_n12, mul_y0y1_n11,
         mul_y0y1_n10, mul_y0y1_n9, mul_y0y1_n8, mul_y0y1_n7, mul_y0y1_n6,
         mul_y0y1_n5, mul_y0y1_n4, mul_y0y1_n3, mul_y0y1_n2, mul_y0y1_n1,
         mul_y0y1_n96, mul_y0y1_n95, mul_y0y1_n94, mul_y0y1_n93, mul_y0y1_n92,
         mul_y0y1_n91, mul_y0y1_n90, mul_y0y1_n89, mul_y0y1_n88, mul_y0y1_n87,
         mul_y0y1_n86, mul_y0y1_n85, mul_y0y1_n84, mul_y0y1_n83, mul_y0y1_n82,
         mul_y0y1_n81, mul_y0y1_n80, mul_y0y1_n79, mul_y0y1_n78, mul_y0y1_n77,
         mul_y0y1_n76, mul_y0y1_n75, mul_y0y1_n74, mul_y0y1_n73, mul_y0y1_n72,
         mul_y0y1_n71, mul_y0y1_n70, mul_y0y1_n69, mul_y0y1_n68, mul_y0y1_n67,
         mul_y0y1_n66, mul_y0y1_n65, mul_y0y1_n64, mul_y0y1_n63, mul_y0y1_n62,
         mul_y0y1_n61, mul_y0y1_n60, mul_y0y1_n59, mul_y0y1_n58, mul_y0y1_n57,
         mul_y0y1_n56, mul_y0y1_n55, mul_y0y1_n54, mul_y0y1_n53, mul_y0y1_n52,
         mul_y0y1_n51, mul_y0y1_n50, mul_y0y1_n49, mul_y0y1_n48, mul_y0y1_n47,
         mul_y0y1_n46, mul_y0y1_n45, mul_y0y1_n44, mul_y0y1_n43, mul_y0y1_n42,
         mul_y0y1_n41, mul_y0y1_n40, mul_y0y1_n39, mul_y0y1_n38, mul_y0y1_n37,
         mul_y0y1_n36, mul_y0y1_n35, mul_y0y1_n34, mul_y0y1_n33,
         mul_y0y1_Xi_mul_Yj_1__0_, mul_y0y1_Xi_mul_Yj_1__1_,
         mul_y0y1_Xi_mul_Yj_1__2_, mul_y0y1_Xi_mul_Yj_1__3_,
         mul_y0y1_Xi_mul_Yj_2__0_, mul_y0y1_Xi_mul_Yj_2__1_,
         mul_y0y1_Xi_mul_Yj_2__2_, mul_y0y1_Xi_mul_Yj_2__3_,
         mul_y0y1_Xi_mul_Yj_3__0_, mul_y0y1_Xi_mul_Yj_3__1_,
         mul_y0y1_Xi_mul_Yj_3__2_, mul_y0y1_Xi_mul_Yj_3__3_,
         mul_y0y1_Xi_mul_Yj_4__0_, mul_y0y1_Xi_mul_Yj_4__1_,
         mul_y0y1_Xi_mul_Yj_4__2_, mul_y0y1_Xi_mul_Yj_4__3_,
         mul_y0y1_Xi_mul_Yj_6__0_, mul_y0y1_Xi_mul_Yj_6__1_,
         mul_y0y1_Xi_mul_Yj_6__2_, mul_y0y1_Xi_mul_Yj_6__3_,
         mul_y0y1_Xi_mul_Yj_7__0_, mul_y0y1_Xi_mul_Yj_7__1_,
         mul_y0y1_Xi_mul_Yj_7__2_, mul_y0y1_Xi_mul_Yj_7__3_,
         mul_y0y1_Xi_mul_Yj_8__0_, mul_y0y1_Xi_mul_Yj_8__1_,
         mul_y0y1_Xi_mul_Yj_8__2_, mul_y0y1_Xi_mul_Yj_8__3_,
         mul_y0y1_Xi_mul_Yj_9__0_, mul_y0y1_Xi_mul_Yj_9__1_,
         mul_y0y1_Xi_mul_Yj_9__2_, mul_y0y1_Xi_mul_Yj_9__3_,
         mul_y0y1_Xi_mul_Yj_11__0_, mul_y0y1_Xi_mul_Yj_11__1_,
         mul_y0y1_Xi_mul_Yj_11__2_, mul_y0y1_Xi_mul_Yj_11__3_,
         mul_y0y1_Xi_mul_Yj_12__0_, mul_y0y1_Xi_mul_Yj_12__1_,
         mul_y0y1_Xi_mul_Yj_12__2_, mul_y0y1_Xi_mul_Yj_12__3_,
         mul_y0y1_Xi_mul_Yj_13__0_, mul_y0y1_Xi_mul_Yj_13__1_,
         mul_y0y1_Xi_mul_Yj_13__2_, mul_y0y1_Xi_mul_Yj_13__3_,
         mul_y0y1_Xi_mul_Yj_14__0_, mul_y0y1_Xi_mul_Yj_14__1_,
         mul_y0y1_Xi_mul_Yj_14__2_, mul_y0y1_Xi_mul_Yj_14__3_,
         mul_y0y1_gf4_mul_3_3_n77, mul_y0y1_gf4_mul_3_3_n76,
         mul_y0y1_gf4_mul_3_3_n75, mul_y0y1_gf4_mul_3_3_n74,
         mul_y0y1_gf4_mul_3_3_n73, mul_y0y1_gf4_mul_3_3_n72,
         mul_y0y1_gf4_mul_3_3_n71, mul_y0y1_gf4_mul_3_3_n70,
         mul_y0y1_gf4_mul_3_3_n69, mul_y0y1_gf4_mul_3_3_n68,
         mul_y0y1_gf4_mul_3_3_n67, mul_y0y1_gf4_mul_3_3_n66,
         mul_y0y1_gf4_mul_3_3_n65, mul_y0y1_gf4_mul_3_3_n64,
         mul_y0y1_gf4_mul_3_3_n63, mul_y0y1_gf4_mul_3_3_n62,
         mul_y0y1_gf4_mul_3_3_n61, mul_y0y1_gf4_mul_3_3_n60,
         mul_y0y1_gf4_mul_3_3_n59, mul_y0y1_gf4_mul_3_3_n58,
         mul_y0y1_gf4_mul_3_3_n57, mul_y0y1_gf4_mul_3_3_n56,
         mul_y0y1_gf4_mul_3_3_n55, mul_y0y1_gf4_mul_3_3_n54,
         mul_y0y1_gf4_mul_3_3_n53, mul_y0y1_gf4_mul_3_2_n77,
         mul_y0y1_gf4_mul_3_2_n76, mul_y0y1_gf4_mul_3_2_n75,
         mul_y0y1_gf4_mul_3_2_n74, mul_y0y1_gf4_mul_3_2_n73,
         mul_y0y1_gf4_mul_3_2_n72, mul_y0y1_gf4_mul_3_2_n71,
         mul_y0y1_gf4_mul_3_2_n70, mul_y0y1_gf4_mul_3_2_n69,
         mul_y0y1_gf4_mul_3_2_n68, mul_y0y1_gf4_mul_3_2_n67,
         mul_y0y1_gf4_mul_3_2_n66, mul_y0y1_gf4_mul_3_2_n65,
         mul_y0y1_gf4_mul_3_2_n64, mul_y0y1_gf4_mul_3_2_n63,
         mul_y0y1_gf4_mul_3_2_n62, mul_y0y1_gf4_mul_3_2_n61,
         mul_y0y1_gf4_mul_3_2_n60, mul_y0y1_gf4_mul_3_2_n59,
         mul_y0y1_gf4_mul_3_2_n58, mul_y0y1_gf4_mul_3_2_n57,
         mul_y0y1_gf4_mul_3_2_n56, mul_y0y1_gf4_mul_3_2_n55,
         mul_y0y1_gf4_mul_3_2_n54, mul_y0y1_gf4_mul_3_2_n53,
         mul_y0y1_gf4_mul_3_1_n77, mul_y0y1_gf4_mul_3_1_n76,
         mul_y0y1_gf4_mul_3_1_n75, mul_y0y1_gf4_mul_3_1_n74,
         mul_y0y1_gf4_mul_3_1_n73, mul_y0y1_gf4_mul_3_1_n72,
         mul_y0y1_gf4_mul_3_1_n71, mul_y0y1_gf4_mul_3_1_n70,
         mul_y0y1_gf4_mul_3_1_n69, mul_y0y1_gf4_mul_3_1_n68,
         mul_y0y1_gf4_mul_3_1_n67, mul_y0y1_gf4_mul_3_1_n66,
         mul_y0y1_gf4_mul_3_1_n65, mul_y0y1_gf4_mul_3_1_n64,
         mul_y0y1_gf4_mul_3_1_n63, mul_y0y1_gf4_mul_3_1_n62,
         mul_y0y1_gf4_mul_3_1_n61, mul_y0y1_gf4_mul_3_1_n60,
         mul_y0y1_gf4_mul_3_1_n59, mul_y0y1_gf4_mul_3_1_n58,
         mul_y0y1_gf4_mul_3_1_n57, mul_y0y1_gf4_mul_3_1_n56,
         mul_y0y1_gf4_mul_3_1_n55, mul_y0y1_gf4_mul_3_1_n54,
         mul_y0y1_gf4_mul_3_1_n53, mul_y0y1_gf4_mul_3_0_n77,
         mul_y0y1_gf4_mul_3_0_n76, mul_y0y1_gf4_mul_3_0_n75,
         mul_y0y1_gf4_mul_3_0_n74, mul_y0y1_gf4_mul_3_0_n73,
         mul_y0y1_gf4_mul_3_0_n72, mul_y0y1_gf4_mul_3_0_n71,
         mul_y0y1_gf4_mul_3_0_n70, mul_y0y1_gf4_mul_3_0_n69,
         mul_y0y1_gf4_mul_3_0_n68, mul_y0y1_gf4_mul_3_0_n67,
         mul_y0y1_gf4_mul_3_0_n66, mul_y0y1_gf4_mul_3_0_n65,
         mul_y0y1_gf4_mul_3_0_n64, mul_y0y1_gf4_mul_3_0_n63,
         mul_y0y1_gf4_mul_3_0_n62, mul_y0y1_gf4_mul_3_0_n61,
         mul_y0y1_gf4_mul_3_0_n60, mul_y0y1_gf4_mul_3_0_n59,
         mul_y0y1_gf4_mul_3_0_n58, mul_y0y1_gf4_mul_3_0_n57,
         mul_y0y1_gf4_mul_3_0_n56, mul_y0y1_gf4_mul_3_0_n55,
         mul_y0y1_gf4_mul_3_0_n54, mul_y0y1_gf4_mul_3_0_n53,
         mul_y0y1_gf4_mul_2_3_n77, mul_y0y1_gf4_mul_2_3_n76,
         mul_y0y1_gf4_mul_2_3_n75, mul_y0y1_gf4_mul_2_3_n74,
         mul_y0y1_gf4_mul_2_3_n73, mul_y0y1_gf4_mul_2_3_n72,
         mul_y0y1_gf4_mul_2_3_n71, mul_y0y1_gf4_mul_2_3_n70,
         mul_y0y1_gf4_mul_2_3_n69, mul_y0y1_gf4_mul_2_3_n68,
         mul_y0y1_gf4_mul_2_3_n67, mul_y0y1_gf4_mul_2_3_n66,
         mul_y0y1_gf4_mul_2_3_n65, mul_y0y1_gf4_mul_2_3_n64,
         mul_y0y1_gf4_mul_2_3_n63, mul_y0y1_gf4_mul_2_3_n62,
         mul_y0y1_gf4_mul_2_3_n61, mul_y0y1_gf4_mul_2_3_n60,
         mul_y0y1_gf4_mul_2_3_n59, mul_y0y1_gf4_mul_2_3_n58,
         mul_y0y1_gf4_mul_2_3_n57, mul_y0y1_gf4_mul_2_3_n56,
         mul_y0y1_gf4_mul_2_3_n55, mul_y0y1_gf4_mul_2_3_n54,
         mul_y0y1_gf4_mul_2_3_n53, mul_y0y1_gf4_mul_2_2_n77,
         mul_y0y1_gf4_mul_2_2_n76, mul_y0y1_gf4_mul_2_2_n75,
         mul_y0y1_gf4_mul_2_2_n74, mul_y0y1_gf4_mul_2_2_n73,
         mul_y0y1_gf4_mul_2_2_n72, mul_y0y1_gf4_mul_2_2_n71,
         mul_y0y1_gf4_mul_2_2_n70, mul_y0y1_gf4_mul_2_2_n69,
         mul_y0y1_gf4_mul_2_2_n68, mul_y0y1_gf4_mul_2_2_n67,
         mul_y0y1_gf4_mul_2_2_n66, mul_y0y1_gf4_mul_2_2_n65,
         mul_y0y1_gf4_mul_2_2_n64, mul_y0y1_gf4_mul_2_2_n63,
         mul_y0y1_gf4_mul_2_2_n62, mul_y0y1_gf4_mul_2_2_n61,
         mul_y0y1_gf4_mul_2_2_n60, mul_y0y1_gf4_mul_2_2_n59,
         mul_y0y1_gf4_mul_2_2_n58, mul_y0y1_gf4_mul_2_2_n57,
         mul_y0y1_gf4_mul_2_2_n56, mul_y0y1_gf4_mul_2_2_n55,
         mul_y0y1_gf4_mul_2_2_n54, mul_y0y1_gf4_mul_2_2_n53,
         mul_y0y1_gf4_mul_2_1_n77, mul_y0y1_gf4_mul_2_1_n76,
         mul_y0y1_gf4_mul_2_1_n75, mul_y0y1_gf4_mul_2_1_n74,
         mul_y0y1_gf4_mul_2_1_n73, mul_y0y1_gf4_mul_2_1_n72,
         mul_y0y1_gf4_mul_2_1_n71, mul_y0y1_gf4_mul_2_1_n70,
         mul_y0y1_gf4_mul_2_1_n69, mul_y0y1_gf4_mul_2_1_n68,
         mul_y0y1_gf4_mul_2_1_n67, mul_y0y1_gf4_mul_2_1_n66,
         mul_y0y1_gf4_mul_2_1_n65, mul_y0y1_gf4_mul_2_1_n64,
         mul_y0y1_gf4_mul_2_1_n63, mul_y0y1_gf4_mul_2_1_n62,
         mul_y0y1_gf4_mul_2_1_n61, mul_y0y1_gf4_mul_2_1_n60,
         mul_y0y1_gf4_mul_2_1_n59, mul_y0y1_gf4_mul_2_1_n58,
         mul_y0y1_gf4_mul_2_1_n57, mul_y0y1_gf4_mul_2_1_n56,
         mul_y0y1_gf4_mul_2_1_n55, mul_y0y1_gf4_mul_2_1_n54,
         mul_y0y1_gf4_mul_2_1_n53, mul_y0y1_gf4_mul_2_0_n77,
         mul_y0y1_gf4_mul_2_0_n76, mul_y0y1_gf4_mul_2_0_n75,
         mul_y0y1_gf4_mul_2_0_n74, mul_y0y1_gf4_mul_2_0_n73,
         mul_y0y1_gf4_mul_2_0_n72, mul_y0y1_gf4_mul_2_0_n71,
         mul_y0y1_gf4_mul_2_0_n70, mul_y0y1_gf4_mul_2_0_n69,
         mul_y0y1_gf4_mul_2_0_n68, mul_y0y1_gf4_mul_2_0_n67,
         mul_y0y1_gf4_mul_2_0_n66, mul_y0y1_gf4_mul_2_0_n65,
         mul_y0y1_gf4_mul_2_0_n64, mul_y0y1_gf4_mul_2_0_n63,
         mul_y0y1_gf4_mul_2_0_n62, mul_y0y1_gf4_mul_2_0_n61,
         mul_y0y1_gf4_mul_2_0_n60, mul_y0y1_gf4_mul_2_0_n59,
         mul_y0y1_gf4_mul_2_0_n58, mul_y0y1_gf4_mul_2_0_n57,
         mul_y0y1_gf4_mul_2_0_n56, mul_y0y1_gf4_mul_2_0_n55,
         mul_y0y1_gf4_mul_2_0_n54, mul_y0y1_gf4_mul_2_0_n53,
         mul_y0y1_gf4_mul_1_3_n77, mul_y0y1_gf4_mul_1_3_n76,
         mul_y0y1_gf4_mul_1_3_n75, mul_y0y1_gf4_mul_1_3_n74,
         mul_y0y1_gf4_mul_1_3_n73, mul_y0y1_gf4_mul_1_3_n72,
         mul_y0y1_gf4_mul_1_3_n71, mul_y0y1_gf4_mul_1_3_n70,
         mul_y0y1_gf4_mul_1_3_n69, mul_y0y1_gf4_mul_1_3_n68,
         mul_y0y1_gf4_mul_1_3_n67, mul_y0y1_gf4_mul_1_3_n66,
         mul_y0y1_gf4_mul_1_3_n65, mul_y0y1_gf4_mul_1_3_n64,
         mul_y0y1_gf4_mul_1_3_n63, mul_y0y1_gf4_mul_1_3_n62,
         mul_y0y1_gf4_mul_1_3_n61, mul_y0y1_gf4_mul_1_3_n60,
         mul_y0y1_gf4_mul_1_3_n59, mul_y0y1_gf4_mul_1_3_n58,
         mul_y0y1_gf4_mul_1_3_n57, mul_y0y1_gf4_mul_1_3_n56,
         mul_y0y1_gf4_mul_1_3_n55, mul_y0y1_gf4_mul_1_3_n54,
         mul_y0y1_gf4_mul_1_3_n53, mul_y0y1_gf4_mul_1_2_n77,
         mul_y0y1_gf4_mul_1_2_n76, mul_y0y1_gf4_mul_1_2_n75,
         mul_y0y1_gf4_mul_1_2_n74, mul_y0y1_gf4_mul_1_2_n73,
         mul_y0y1_gf4_mul_1_2_n72, mul_y0y1_gf4_mul_1_2_n71,
         mul_y0y1_gf4_mul_1_2_n70, mul_y0y1_gf4_mul_1_2_n69,
         mul_y0y1_gf4_mul_1_2_n68, mul_y0y1_gf4_mul_1_2_n67,
         mul_y0y1_gf4_mul_1_2_n66, mul_y0y1_gf4_mul_1_2_n65,
         mul_y0y1_gf4_mul_1_2_n64, mul_y0y1_gf4_mul_1_2_n63,
         mul_y0y1_gf4_mul_1_2_n62, mul_y0y1_gf4_mul_1_2_n61,
         mul_y0y1_gf4_mul_1_2_n60, mul_y0y1_gf4_mul_1_2_n59,
         mul_y0y1_gf4_mul_1_2_n58, mul_y0y1_gf4_mul_1_2_n57,
         mul_y0y1_gf4_mul_1_2_n56, mul_y0y1_gf4_mul_1_2_n55,
         mul_y0y1_gf4_mul_1_2_n54, mul_y0y1_gf4_mul_1_2_n53,
         mul_y0y1_gf4_mul_1_1_n77, mul_y0y1_gf4_mul_1_1_n76,
         mul_y0y1_gf4_mul_1_1_n75, mul_y0y1_gf4_mul_1_1_n74,
         mul_y0y1_gf4_mul_1_1_n73, mul_y0y1_gf4_mul_1_1_n72,
         mul_y0y1_gf4_mul_1_1_n71, mul_y0y1_gf4_mul_1_1_n70,
         mul_y0y1_gf4_mul_1_1_n69, mul_y0y1_gf4_mul_1_1_n68,
         mul_y0y1_gf4_mul_1_1_n67, mul_y0y1_gf4_mul_1_1_n66,
         mul_y0y1_gf4_mul_1_1_n65, mul_y0y1_gf4_mul_1_1_n64,
         mul_y0y1_gf4_mul_1_1_n63, mul_y0y1_gf4_mul_1_1_n62,
         mul_y0y1_gf4_mul_1_1_n61, mul_y0y1_gf4_mul_1_1_n60,
         mul_y0y1_gf4_mul_1_1_n59, mul_y0y1_gf4_mul_1_1_n58,
         mul_y0y1_gf4_mul_1_1_n57, mul_y0y1_gf4_mul_1_1_n56,
         mul_y0y1_gf4_mul_1_1_n55, mul_y0y1_gf4_mul_1_1_n54,
         mul_y0y1_gf4_mul_1_1_n53, mul_y0y1_gf4_mul_1_0_n77,
         mul_y0y1_gf4_mul_1_0_n76, mul_y0y1_gf4_mul_1_0_n75,
         mul_y0y1_gf4_mul_1_0_n74, mul_y0y1_gf4_mul_1_0_n73,
         mul_y0y1_gf4_mul_1_0_n72, mul_y0y1_gf4_mul_1_0_n71,
         mul_y0y1_gf4_mul_1_0_n70, mul_y0y1_gf4_mul_1_0_n69,
         mul_y0y1_gf4_mul_1_0_n68, mul_y0y1_gf4_mul_1_0_n67,
         mul_y0y1_gf4_mul_1_0_n66, mul_y0y1_gf4_mul_1_0_n65,
         mul_y0y1_gf4_mul_1_0_n64, mul_y0y1_gf4_mul_1_0_n63,
         mul_y0y1_gf4_mul_1_0_n62, mul_y0y1_gf4_mul_1_0_n61,
         mul_y0y1_gf4_mul_1_0_n60, mul_y0y1_gf4_mul_1_0_n59,
         mul_y0y1_gf4_mul_1_0_n58, mul_y0y1_gf4_mul_1_0_n57,
         mul_y0y1_gf4_mul_1_0_n56, mul_y0y1_gf4_mul_1_0_n55,
         mul_y0y1_gf4_mul_1_0_n54, mul_y0y1_gf4_mul_1_0_n53,
         mul_y0y1_gf4_mul_0_3_n77, mul_y0y1_gf4_mul_0_3_n76,
         mul_y0y1_gf4_mul_0_3_n75, mul_y0y1_gf4_mul_0_3_n74,
         mul_y0y1_gf4_mul_0_3_n73, mul_y0y1_gf4_mul_0_3_n72,
         mul_y0y1_gf4_mul_0_3_n71, mul_y0y1_gf4_mul_0_3_n70,
         mul_y0y1_gf4_mul_0_3_n69, mul_y0y1_gf4_mul_0_3_n68,
         mul_y0y1_gf4_mul_0_3_n67, mul_y0y1_gf4_mul_0_3_n66,
         mul_y0y1_gf4_mul_0_3_n65, mul_y0y1_gf4_mul_0_3_n64,
         mul_y0y1_gf4_mul_0_3_n63, mul_y0y1_gf4_mul_0_3_n62,
         mul_y0y1_gf4_mul_0_3_n61, mul_y0y1_gf4_mul_0_3_n60,
         mul_y0y1_gf4_mul_0_3_n59, mul_y0y1_gf4_mul_0_3_n58,
         mul_y0y1_gf4_mul_0_3_n57, mul_y0y1_gf4_mul_0_3_n56,
         mul_y0y1_gf4_mul_0_3_n55, mul_y0y1_gf4_mul_0_3_n54,
         mul_y0y1_gf4_mul_0_3_n53, mul_y0y1_gf4_mul_0_2_n77,
         mul_y0y1_gf4_mul_0_2_n76, mul_y0y1_gf4_mul_0_2_n75,
         mul_y0y1_gf4_mul_0_2_n74, mul_y0y1_gf4_mul_0_2_n73,
         mul_y0y1_gf4_mul_0_2_n72, mul_y0y1_gf4_mul_0_2_n71,
         mul_y0y1_gf4_mul_0_2_n70, mul_y0y1_gf4_mul_0_2_n69,
         mul_y0y1_gf4_mul_0_2_n68, mul_y0y1_gf4_mul_0_2_n67,
         mul_y0y1_gf4_mul_0_2_n66, mul_y0y1_gf4_mul_0_2_n65,
         mul_y0y1_gf4_mul_0_2_n64, mul_y0y1_gf4_mul_0_2_n63,
         mul_y0y1_gf4_mul_0_2_n62, mul_y0y1_gf4_mul_0_2_n61,
         mul_y0y1_gf4_mul_0_2_n60, mul_y0y1_gf4_mul_0_2_n59,
         mul_y0y1_gf4_mul_0_2_n58, mul_y0y1_gf4_mul_0_2_n57,
         mul_y0y1_gf4_mul_0_2_n56, mul_y0y1_gf4_mul_0_2_n55,
         mul_y0y1_gf4_mul_0_2_n54, mul_y0y1_gf4_mul_0_2_n53,
         mul_y0y1_gf4_mul_0_1_n77, mul_y0y1_gf4_mul_0_1_n76,
         mul_y0y1_gf4_mul_0_1_n75, mul_y0y1_gf4_mul_0_1_n74,
         mul_y0y1_gf4_mul_0_1_n73, mul_y0y1_gf4_mul_0_1_n72,
         mul_y0y1_gf4_mul_0_1_n71, mul_y0y1_gf4_mul_0_1_n70,
         mul_y0y1_gf4_mul_0_1_n69, mul_y0y1_gf4_mul_0_1_n68,
         mul_y0y1_gf4_mul_0_1_n67, mul_y0y1_gf4_mul_0_1_n66,
         mul_y0y1_gf4_mul_0_1_n65, mul_y0y1_gf4_mul_0_1_n64,
         mul_y0y1_gf4_mul_0_1_n63, mul_y0y1_gf4_mul_0_1_n62,
         mul_y0y1_gf4_mul_0_1_n61, mul_y0y1_gf4_mul_0_1_n60,
         mul_y0y1_gf4_mul_0_1_n59, mul_y0y1_gf4_mul_0_1_n58,
         mul_y0y1_gf4_mul_0_1_n57, mul_y0y1_gf4_mul_0_1_n56,
         mul_y0y1_gf4_mul_0_1_n55, mul_y0y1_gf4_mul_0_1_n54,
         mul_y0y1_gf4_mul_0_1_n53, mul_y0y1_gf4_mul_0_0_n77,
         mul_y0y1_gf4_mul_0_0_n76, mul_y0y1_gf4_mul_0_0_n75,
         mul_y0y1_gf4_mul_0_0_n74, mul_y0y1_gf4_mul_0_0_n73,
         mul_y0y1_gf4_mul_0_0_n72, mul_y0y1_gf4_mul_0_0_n71,
         mul_y0y1_gf4_mul_0_0_n70, mul_y0y1_gf4_mul_0_0_n69,
         mul_y0y1_gf4_mul_0_0_n68, mul_y0y1_gf4_mul_0_0_n67,
         mul_y0y1_gf4_mul_0_0_n66, mul_y0y1_gf4_mul_0_0_n65,
         mul_y0y1_gf4_mul_0_0_n64, mul_y0y1_gf4_mul_0_0_n63,
         mul_y0y1_gf4_mul_0_0_n62, mul_y0y1_gf4_mul_0_0_n61,
         mul_y0y1_gf4_mul_0_0_n60, mul_y0y1_gf4_mul_0_0_n59,
         mul_y0y1_gf4_mul_0_0_n58, mul_y0y1_gf4_mul_0_0_n57,
         mul_y0y1_gf4_mul_0_0_n56, mul_y0y1_gf4_mul_0_0_n55,
         mul_y0y1_gf4_mul_0_0_n54, mul_y0y1_gf4_mul_0_0_n53, inverter_gf24_n4,
         inverter_gf24_n3, inverter_gf24_n2, inverter_gf24_n1,
         inverter_gf24_n16, inverter_gf24_n15, inverter_gf24_n14,
         inverter_gf24_n13, inverter_gf24_n12, inverter_gf24_n11,
         inverter_gf24_n10, inverter_gf24_n9, inverter_gf24_n8,
         inverter_gf24_n7, inverter_gf24_n6, inverter_gf24_n5,
         inverter_gf24_d_0__0_, inverter_gf24_d_1__0_, inverter_gf24_d_2__0_,
         inverter_gf24_d_3__0_, inverter_gf24_ExDP_0__0_,
         inverter_gf24_ExDP_0__1_, inverter_gf24_ExDP_1__0_,
         inverter_gf24_ExDP_1__1_, inverter_gf24_ExDP_2__0_,
         inverter_gf24_ExDP_2__1_, inverter_gf24_ExDP_3__0_,
         inverter_gf24_ExDP_3__1_, inverter_gf24_a_mul_b_n16,
         inverter_gf24_a_mul_b_n15, inverter_gf24_a_mul_b_n14,
         inverter_gf24_a_mul_b_n13, inverter_gf24_a_mul_b_n12,
         inverter_gf24_a_mul_b_n11, inverter_gf24_a_mul_b_n10,
         inverter_gf24_a_mul_b_n9, inverter_gf24_a_mul_b_n8,
         inverter_gf24_a_mul_b_n7, inverter_gf24_a_mul_b_n6,
         inverter_gf24_a_mul_b_n5, inverter_gf24_a_mul_b_n4,
         inverter_gf24_a_mul_b_n3, inverter_gf24_a_mul_b_n2,
         inverter_gf24_a_mul_b_n1, inverter_gf24_a_mul_b_n48,
         inverter_gf24_a_mul_b_n47, inverter_gf24_a_mul_b_n46,
         inverter_gf24_a_mul_b_n45, inverter_gf24_a_mul_b_n44,
         inverter_gf24_a_mul_b_n43, inverter_gf24_a_mul_b_n42,
         inverter_gf24_a_mul_b_n41, inverter_gf24_a_mul_b_n40,
         inverter_gf24_a_mul_b_n39, inverter_gf24_a_mul_b_n38,
         inverter_gf24_a_mul_b_n37, inverter_gf24_a_mul_b_n36,
         inverter_gf24_a_mul_b_n35, inverter_gf24_a_mul_b_n34,
         inverter_gf24_a_mul_b_n33, inverter_gf24_a_mul_b_n32,
         inverter_gf24_a_mul_b_n31, inverter_gf24_a_mul_b_n30,
         inverter_gf24_a_mul_b_n29, inverter_gf24_a_mul_b_n28,
         inverter_gf24_a_mul_b_n27, inverter_gf24_a_mul_b_n26,
         inverter_gf24_a_mul_b_n25, inverter_gf24_a_mul_b_n24,
         inverter_gf24_a_mul_b_n23, inverter_gf24_a_mul_b_n22,
         inverter_gf24_a_mul_b_n21, inverter_gf24_a_mul_b_n20,
         inverter_gf24_a_mul_b_n19, inverter_gf24_a_mul_b_n18,
         inverter_gf24_a_mul_b_n17, inverter_gf24_a_mul_b_Xi_mul_Yj_1__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_1__1_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_2__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_2__1_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_3__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_3__1_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_4__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_4__1_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_6__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_6__1_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_7__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_7__1_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_8__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_8__1_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_9__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_9__1_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_11__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_11__1_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_12__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_12__1_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_13__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_13__1_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_14__0_,
         inverter_gf24_a_mul_b_Xi_mul_Yj_14__1_,
         inverter_gf24_a_mul_b_gf2_mul_3_3_n15,
         inverter_gf24_a_mul_b_gf2_mul_3_3_n14,
         inverter_gf24_a_mul_b_gf2_mul_3_3_n13,
         inverter_gf24_a_mul_b_gf2_mul_3_3_n12,
         inverter_gf24_a_mul_b_gf2_mul_3_3_n11,
         inverter_gf24_a_mul_b_gf2_mul_3_2_n15,
         inverter_gf24_a_mul_b_gf2_mul_3_2_n14,
         inverter_gf24_a_mul_b_gf2_mul_3_2_n13,
         inverter_gf24_a_mul_b_gf2_mul_3_2_n12,
         inverter_gf24_a_mul_b_gf2_mul_3_2_n11,
         inverter_gf24_a_mul_b_gf2_mul_3_1_n15,
         inverter_gf24_a_mul_b_gf2_mul_3_1_n14,
         inverter_gf24_a_mul_b_gf2_mul_3_1_n13,
         inverter_gf24_a_mul_b_gf2_mul_3_1_n12,
         inverter_gf24_a_mul_b_gf2_mul_3_1_n11,
         inverter_gf24_a_mul_b_gf2_mul_3_0_n15,
         inverter_gf24_a_mul_b_gf2_mul_3_0_n14,
         inverter_gf24_a_mul_b_gf2_mul_3_0_n13,
         inverter_gf24_a_mul_b_gf2_mul_3_0_n12,
         inverter_gf24_a_mul_b_gf2_mul_3_0_n11,
         inverter_gf24_a_mul_b_gf2_mul_2_3_n15,
         inverter_gf24_a_mul_b_gf2_mul_2_3_n14,
         inverter_gf24_a_mul_b_gf2_mul_2_3_n13,
         inverter_gf24_a_mul_b_gf2_mul_2_3_n12,
         inverter_gf24_a_mul_b_gf2_mul_2_3_n11,
         inverter_gf24_a_mul_b_gf2_mul_2_2_n15,
         inverter_gf24_a_mul_b_gf2_mul_2_2_n14,
         inverter_gf24_a_mul_b_gf2_mul_2_2_n13,
         inverter_gf24_a_mul_b_gf2_mul_2_2_n12,
         inverter_gf24_a_mul_b_gf2_mul_2_2_n11,
         inverter_gf24_a_mul_b_gf2_mul_2_1_n15,
         inverter_gf24_a_mul_b_gf2_mul_2_1_n14,
         inverter_gf24_a_mul_b_gf2_mul_2_1_n13,
         inverter_gf24_a_mul_b_gf2_mul_2_1_n12,
         inverter_gf24_a_mul_b_gf2_mul_2_1_n11,
         inverter_gf24_a_mul_b_gf2_mul_2_0_n15,
         inverter_gf24_a_mul_b_gf2_mul_2_0_n14,
         inverter_gf24_a_mul_b_gf2_mul_2_0_n13,
         inverter_gf24_a_mul_b_gf2_mul_2_0_n12,
         inverter_gf24_a_mul_b_gf2_mul_2_0_n11,
         inverter_gf24_a_mul_b_gf2_mul_1_3_n15,
         inverter_gf24_a_mul_b_gf2_mul_1_3_n14,
         inverter_gf24_a_mul_b_gf2_mul_1_3_n13,
         inverter_gf24_a_mul_b_gf2_mul_1_3_n12,
         inverter_gf24_a_mul_b_gf2_mul_1_3_n11,
         inverter_gf24_a_mul_b_gf2_mul_1_2_n15,
         inverter_gf24_a_mul_b_gf2_mul_1_2_n14,
         inverter_gf24_a_mul_b_gf2_mul_1_2_n13,
         inverter_gf24_a_mul_b_gf2_mul_1_2_n12,
         inverter_gf24_a_mul_b_gf2_mul_1_2_n11,
         inverter_gf24_a_mul_b_gf2_mul_1_1_n15,
         inverter_gf24_a_mul_b_gf2_mul_1_1_n14,
         inverter_gf24_a_mul_b_gf2_mul_1_1_n13,
         inverter_gf24_a_mul_b_gf2_mul_1_1_n12,
         inverter_gf24_a_mul_b_gf2_mul_1_1_n11,
         inverter_gf24_a_mul_b_gf2_mul_1_0_n15,
         inverter_gf24_a_mul_b_gf2_mul_1_0_n14,
         inverter_gf24_a_mul_b_gf2_mul_1_0_n13,
         inverter_gf24_a_mul_b_gf2_mul_1_0_n12,
         inverter_gf24_a_mul_b_gf2_mul_1_0_n11,
         inverter_gf24_a_mul_b_gf2_mul_0_3_n15,
         inverter_gf24_a_mul_b_gf2_mul_0_3_n14,
         inverter_gf24_a_mul_b_gf2_mul_0_3_n13,
         inverter_gf24_a_mul_b_gf2_mul_0_3_n12,
         inverter_gf24_a_mul_b_gf2_mul_0_3_n11,
         inverter_gf24_a_mul_b_gf2_mul_0_2_n15,
         inverter_gf24_a_mul_b_gf2_mul_0_2_n14,
         inverter_gf24_a_mul_b_gf2_mul_0_2_n13,
         inverter_gf24_a_mul_b_gf2_mul_0_2_n12,
         inverter_gf24_a_mul_b_gf2_mul_0_2_n11,
         inverter_gf24_a_mul_b_gf2_mul_0_1_n15,
         inverter_gf24_a_mul_b_gf2_mul_0_1_n14,
         inverter_gf24_a_mul_b_gf2_mul_0_1_n13,
         inverter_gf24_a_mul_b_gf2_mul_0_1_n12,
         inverter_gf24_a_mul_b_gf2_mul_0_1_n11,
         inverter_gf24_a_mul_b_gf2_mul_0_0_n15,
         inverter_gf24_a_mul_b_gf2_mul_0_0_n14,
         inverter_gf24_a_mul_b_gf2_mul_0_0_n13,
         inverter_gf24_a_mul_b_gf2_mul_0_0_n12,
         inverter_gf24_a_mul_b_gf2_mul_0_0_n11, inverter_gf24_a_mul_e_n64,
         inverter_gf24_a_mul_e_n63, inverter_gf24_a_mul_e_n62,
         inverter_gf24_a_mul_e_n61, inverter_gf24_a_mul_e_n60,
         inverter_gf24_a_mul_e_n59, inverter_gf24_a_mul_e_n58,
         inverter_gf24_a_mul_e_n57, inverter_gf24_a_mul_e_n56,
         inverter_gf24_a_mul_e_n55, inverter_gf24_a_mul_e_n54,
         inverter_gf24_a_mul_e_n53, inverter_gf24_a_mul_e_n52,
         inverter_gf24_a_mul_e_n51, inverter_gf24_a_mul_e_n50,
         inverter_gf24_a_mul_e_n49, inverter_gf24_a_mul_e_n48,
         inverter_gf24_a_mul_e_n47, inverter_gf24_a_mul_e_n46,
         inverter_gf24_a_mul_e_n45, inverter_gf24_a_mul_e_n44,
         inverter_gf24_a_mul_e_n43, inverter_gf24_a_mul_e_n42,
         inverter_gf24_a_mul_e_n41, inverter_gf24_a_mul_e_n40,
         inverter_gf24_a_mul_e_n39, inverter_gf24_a_mul_e_n38,
         inverter_gf24_a_mul_e_n37, inverter_gf24_a_mul_e_n36,
         inverter_gf24_a_mul_e_n35, inverter_gf24_a_mul_e_n34,
         inverter_gf24_a_mul_e_n33, inverter_gf24_a_mul_e_n32,
         inverter_gf24_a_mul_e_n31, inverter_gf24_a_mul_e_n30,
         inverter_gf24_a_mul_e_n29, inverter_gf24_a_mul_e_n28,
         inverter_gf24_a_mul_e_n27, inverter_gf24_a_mul_e_n26,
         inverter_gf24_a_mul_e_n25, inverter_gf24_a_mul_e_n24,
         inverter_gf24_a_mul_e_n23, inverter_gf24_a_mul_e_n22,
         inverter_gf24_a_mul_e_n21, inverter_gf24_a_mul_e_n20,
         inverter_gf24_a_mul_e_n19, inverter_gf24_a_mul_e_n18,
         inverter_gf24_a_mul_e_n17, inverter_gf24_a_mul_e_Xi_mul_Yj_1__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_1__1_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_2__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_2__1_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_3__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_3__1_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_4__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_4__1_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_6__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_6__1_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_7__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_7__1_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_8__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_8__1_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_9__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_9__1_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_11__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_11__1_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_12__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_12__1_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_13__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_13__1_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_14__0_,
         inverter_gf24_a_mul_e_Xi_mul_Yj_14__1_,
         inverter_gf24_a_mul_e_gf2_mul_3_3_n15,
         inverter_gf24_a_mul_e_gf2_mul_3_3_n14,
         inverter_gf24_a_mul_e_gf2_mul_3_3_n13,
         inverter_gf24_a_mul_e_gf2_mul_3_3_n12,
         inverter_gf24_a_mul_e_gf2_mul_3_3_n11,
         inverter_gf24_a_mul_e_gf2_mul_3_2_n15,
         inverter_gf24_a_mul_e_gf2_mul_3_2_n14,
         inverter_gf24_a_mul_e_gf2_mul_3_2_n13,
         inverter_gf24_a_mul_e_gf2_mul_3_2_n12,
         inverter_gf24_a_mul_e_gf2_mul_3_2_n11,
         inverter_gf24_a_mul_e_gf2_mul_3_1_n15,
         inverter_gf24_a_mul_e_gf2_mul_3_1_n14,
         inverter_gf24_a_mul_e_gf2_mul_3_1_n13,
         inverter_gf24_a_mul_e_gf2_mul_3_1_n12,
         inverter_gf24_a_mul_e_gf2_mul_3_1_n11,
         inverter_gf24_a_mul_e_gf2_mul_3_0_n15,
         inverter_gf24_a_mul_e_gf2_mul_3_0_n14,
         inverter_gf24_a_mul_e_gf2_mul_3_0_n13,
         inverter_gf24_a_mul_e_gf2_mul_3_0_n12,
         inverter_gf24_a_mul_e_gf2_mul_3_0_n11,
         inverter_gf24_a_mul_e_gf2_mul_2_3_n15,
         inverter_gf24_a_mul_e_gf2_mul_2_3_n14,
         inverter_gf24_a_mul_e_gf2_mul_2_3_n13,
         inverter_gf24_a_mul_e_gf2_mul_2_3_n12,
         inverter_gf24_a_mul_e_gf2_mul_2_3_n11,
         inverter_gf24_a_mul_e_gf2_mul_2_2_n15,
         inverter_gf24_a_mul_e_gf2_mul_2_2_n14,
         inverter_gf24_a_mul_e_gf2_mul_2_2_n13,
         inverter_gf24_a_mul_e_gf2_mul_2_2_n12,
         inverter_gf24_a_mul_e_gf2_mul_2_2_n11,
         inverter_gf24_a_mul_e_gf2_mul_2_1_n15,
         inverter_gf24_a_mul_e_gf2_mul_2_1_n14,
         inverter_gf24_a_mul_e_gf2_mul_2_1_n13,
         inverter_gf24_a_mul_e_gf2_mul_2_1_n12,
         inverter_gf24_a_mul_e_gf2_mul_2_1_n11,
         inverter_gf24_a_mul_e_gf2_mul_2_0_n15,
         inverter_gf24_a_mul_e_gf2_mul_2_0_n14,
         inverter_gf24_a_mul_e_gf2_mul_2_0_n13,
         inverter_gf24_a_mul_e_gf2_mul_2_0_n12,
         inverter_gf24_a_mul_e_gf2_mul_2_0_n11,
         inverter_gf24_a_mul_e_gf2_mul_1_3_n15,
         inverter_gf24_a_mul_e_gf2_mul_1_3_n14,
         inverter_gf24_a_mul_e_gf2_mul_1_3_n13,
         inverter_gf24_a_mul_e_gf2_mul_1_3_n12,
         inverter_gf24_a_mul_e_gf2_mul_1_3_n11,
         inverter_gf24_a_mul_e_gf2_mul_1_2_n15,
         inverter_gf24_a_mul_e_gf2_mul_1_2_n14,
         inverter_gf24_a_mul_e_gf2_mul_1_2_n13,
         inverter_gf24_a_mul_e_gf2_mul_1_2_n12,
         inverter_gf24_a_mul_e_gf2_mul_1_2_n11,
         inverter_gf24_a_mul_e_gf2_mul_1_1_n15,
         inverter_gf24_a_mul_e_gf2_mul_1_1_n14,
         inverter_gf24_a_mul_e_gf2_mul_1_1_n13,
         inverter_gf24_a_mul_e_gf2_mul_1_1_n12,
         inverter_gf24_a_mul_e_gf2_mul_1_1_n11,
         inverter_gf24_a_mul_e_gf2_mul_1_0_n15,
         inverter_gf24_a_mul_e_gf2_mul_1_0_n14,
         inverter_gf24_a_mul_e_gf2_mul_1_0_n13,
         inverter_gf24_a_mul_e_gf2_mul_1_0_n12,
         inverter_gf24_a_mul_e_gf2_mul_1_0_n11,
         inverter_gf24_a_mul_e_gf2_mul_0_3_n15,
         inverter_gf24_a_mul_e_gf2_mul_0_3_n14,
         inverter_gf24_a_mul_e_gf2_mul_0_3_n13,
         inverter_gf24_a_mul_e_gf2_mul_0_3_n12,
         inverter_gf24_a_mul_e_gf2_mul_0_3_n11,
         inverter_gf24_a_mul_e_gf2_mul_0_2_n15,
         inverter_gf24_a_mul_e_gf2_mul_0_2_n14,
         inverter_gf24_a_mul_e_gf2_mul_0_2_n13,
         inverter_gf24_a_mul_e_gf2_mul_0_2_n12,
         inverter_gf24_a_mul_e_gf2_mul_0_2_n11,
         inverter_gf24_a_mul_e_gf2_mul_0_1_n15,
         inverter_gf24_a_mul_e_gf2_mul_0_1_n14,
         inverter_gf24_a_mul_e_gf2_mul_0_1_n13,
         inverter_gf24_a_mul_e_gf2_mul_0_1_n12,
         inverter_gf24_a_mul_e_gf2_mul_0_1_n11,
         inverter_gf24_a_mul_e_gf2_mul_0_0_n15,
         inverter_gf24_a_mul_e_gf2_mul_0_0_n14,
         inverter_gf24_a_mul_e_gf2_mul_0_0_n13,
         inverter_gf24_a_mul_e_gf2_mul_0_0_n12,
         inverter_gf24_a_mul_e_gf2_mul_0_0_n11, inverter_gf24_b_mul_e_n64,
         inverter_gf24_b_mul_e_n63, inverter_gf24_b_mul_e_n62,
         inverter_gf24_b_mul_e_n61, inverter_gf24_b_mul_e_n60,
         inverter_gf24_b_mul_e_n59, inverter_gf24_b_mul_e_n58,
         inverter_gf24_b_mul_e_n57, inverter_gf24_b_mul_e_n56,
         inverter_gf24_b_mul_e_n55, inverter_gf24_b_mul_e_n54,
         inverter_gf24_b_mul_e_n53, inverter_gf24_b_mul_e_n52,
         inverter_gf24_b_mul_e_n51, inverter_gf24_b_mul_e_n50,
         inverter_gf24_b_mul_e_n49, inverter_gf24_b_mul_e_n48,
         inverter_gf24_b_mul_e_n47, inverter_gf24_b_mul_e_n46,
         inverter_gf24_b_mul_e_n45, inverter_gf24_b_mul_e_n44,
         inverter_gf24_b_mul_e_n43, inverter_gf24_b_mul_e_n42,
         inverter_gf24_b_mul_e_n41, inverter_gf24_b_mul_e_n40,
         inverter_gf24_b_mul_e_n39, inverter_gf24_b_mul_e_n38,
         inverter_gf24_b_mul_e_n37, inverter_gf24_b_mul_e_n36,
         inverter_gf24_b_mul_e_n35, inverter_gf24_b_mul_e_n34,
         inverter_gf24_b_mul_e_n33, inverter_gf24_b_mul_e_n32,
         inverter_gf24_b_mul_e_n31, inverter_gf24_b_mul_e_n30,
         inverter_gf24_b_mul_e_n29, inverter_gf24_b_mul_e_n28,
         inverter_gf24_b_mul_e_n27, inverter_gf24_b_mul_e_n26,
         inverter_gf24_b_mul_e_n25, inverter_gf24_b_mul_e_n24,
         inverter_gf24_b_mul_e_n23, inverter_gf24_b_mul_e_n22,
         inverter_gf24_b_mul_e_n21, inverter_gf24_b_mul_e_n20,
         inverter_gf24_b_mul_e_n19, inverter_gf24_b_mul_e_n18,
         inverter_gf24_b_mul_e_n17, inverter_gf24_b_mul_e_Xi_mul_Yj_1__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_1__1_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_2__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_2__1_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_3__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_3__1_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_4__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_4__1_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_6__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_6__1_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_7__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_7__1_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_8__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_8__1_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_9__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_9__1_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_11__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_11__1_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_12__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_12__1_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_13__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_13__1_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_14__0_,
         inverter_gf24_b_mul_e_Xi_mul_Yj_14__1_,
         inverter_gf24_b_mul_e_gf2_mul_3_3_n15,
         inverter_gf24_b_mul_e_gf2_mul_3_3_n14,
         inverter_gf24_b_mul_e_gf2_mul_3_3_n13,
         inverter_gf24_b_mul_e_gf2_mul_3_3_n12,
         inverter_gf24_b_mul_e_gf2_mul_3_3_n11,
         inverter_gf24_b_mul_e_gf2_mul_3_2_n15,
         inverter_gf24_b_mul_e_gf2_mul_3_2_n14,
         inverter_gf24_b_mul_e_gf2_mul_3_2_n13,
         inverter_gf24_b_mul_e_gf2_mul_3_2_n12,
         inverter_gf24_b_mul_e_gf2_mul_3_2_n11,
         inverter_gf24_b_mul_e_gf2_mul_3_1_n15,
         inverter_gf24_b_mul_e_gf2_mul_3_1_n14,
         inverter_gf24_b_mul_e_gf2_mul_3_1_n13,
         inverter_gf24_b_mul_e_gf2_mul_3_1_n12,
         inverter_gf24_b_mul_e_gf2_mul_3_1_n11,
         inverter_gf24_b_mul_e_gf2_mul_3_0_n15,
         inverter_gf24_b_mul_e_gf2_mul_3_0_n14,
         inverter_gf24_b_mul_e_gf2_mul_3_0_n13,
         inverter_gf24_b_mul_e_gf2_mul_3_0_n12,
         inverter_gf24_b_mul_e_gf2_mul_3_0_n11,
         inverter_gf24_b_mul_e_gf2_mul_2_3_n15,
         inverter_gf24_b_mul_e_gf2_mul_2_3_n14,
         inverter_gf24_b_mul_e_gf2_mul_2_3_n13,
         inverter_gf24_b_mul_e_gf2_mul_2_3_n12,
         inverter_gf24_b_mul_e_gf2_mul_2_3_n11,
         inverter_gf24_b_mul_e_gf2_mul_2_2_n15,
         inverter_gf24_b_mul_e_gf2_mul_2_2_n14,
         inverter_gf24_b_mul_e_gf2_mul_2_2_n13,
         inverter_gf24_b_mul_e_gf2_mul_2_2_n12,
         inverter_gf24_b_mul_e_gf2_mul_2_2_n11,
         inverter_gf24_b_mul_e_gf2_mul_2_1_n15,
         inverter_gf24_b_mul_e_gf2_mul_2_1_n14,
         inverter_gf24_b_mul_e_gf2_mul_2_1_n13,
         inverter_gf24_b_mul_e_gf2_mul_2_1_n12,
         inverter_gf24_b_mul_e_gf2_mul_2_1_n11,
         inverter_gf24_b_mul_e_gf2_mul_2_0_n15,
         inverter_gf24_b_mul_e_gf2_mul_2_0_n14,
         inverter_gf24_b_mul_e_gf2_mul_2_0_n13,
         inverter_gf24_b_mul_e_gf2_mul_2_0_n12,
         inverter_gf24_b_mul_e_gf2_mul_2_0_n11,
         inverter_gf24_b_mul_e_gf2_mul_1_3_n15,
         inverter_gf24_b_mul_e_gf2_mul_1_3_n14,
         inverter_gf24_b_mul_e_gf2_mul_1_3_n13,
         inverter_gf24_b_mul_e_gf2_mul_1_3_n12,
         inverter_gf24_b_mul_e_gf2_mul_1_3_n11,
         inverter_gf24_b_mul_e_gf2_mul_1_2_n15,
         inverter_gf24_b_mul_e_gf2_mul_1_2_n14,
         inverter_gf24_b_mul_e_gf2_mul_1_2_n13,
         inverter_gf24_b_mul_e_gf2_mul_1_2_n12,
         inverter_gf24_b_mul_e_gf2_mul_1_2_n11,
         inverter_gf24_b_mul_e_gf2_mul_1_1_n15,
         inverter_gf24_b_mul_e_gf2_mul_1_1_n14,
         inverter_gf24_b_mul_e_gf2_mul_1_1_n13,
         inverter_gf24_b_mul_e_gf2_mul_1_1_n12,
         inverter_gf24_b_mul_e_gf2_mul_1_1_n11,
         inverter_gf24_b_mul_e_gf2_mul_1_0_n15,
         inverter_gf24_b_mul_e_gf2_mul_1_0_n14,
         inverter_gf24_b_mul_e_gf2_mul_1_0_n13,
         inverter_gf24_b_mul_e_gf2_mul_1_0_n12,
         inverter_gf24_b_mul_e_gf2_mul_1_0_n11,
         inverter_gf24_b_mul_e_gf2_mul_0_3_n15,
         inverter_gf24_b_mul_e_gf2_mul_0_3_n14,
         inverter_gf24_b_mul_e_gf2_mul_0_3_n13,
         inverter_gf24_b_mul_e_gf2_mul_0_3_n12,
         inverter_gf24_b_mul_e_gf2_mul_0_3_n11,
         inverter_gf24_b_mul_e_gf2_mul_0_2_n15,
         inverter_gf24_b_mul_e_gf2_mul_0_2_n14,
         inverter_gf24_b_mul_e_gf2_mul_0_2_n13,
         inverter_gf24_b_mul_e_gf2_mul_0_2_n12,
         inverter_gf24_b_mul_e_gf2_mul_0_2_n11,
         inverter_gf24_b_mul_e_gf2_mul_0_1_n15,
         inverter_gf24_b_mul_e_gf2_mul_0_1_n14,
         inverter_gf24_b_mul_e_gf2_mul_0_1_n13,
         inverter_gf24_b_mul_e_gf2_mul_0_1_n12,
         inverter_gf24_b_mul_e_gf2_mul_0_1_n11,
         inverter_gf24_b_mul_e_gf2_mul_0_0_n15,
         inverter_gf24_b_mul_e_gf2_mul_0_0_n14,
         inverter_gf24_b_mul_e_gf2_mul_0_0_n13,
         inverter_gf24_b_mul_e_gf2_mul_0_0_n12,
         inverter_gf24_b_mul_e_gf2_mul_0_0_n11, mult_msb_n128, mult_msb_n127,
         mult_msb_n126, mult_msb_n125, mult_msb_n124, mult_msb_n123,
         mult_msb_n122, mult_msb_n121, mult_msb_n120, mult_msb_n119,
         mult_msb_n118, mult_msb_n117, mult_msb_n116, mult_msb_n115,
         mult_msb_n114, mult_msb_n113, mult_msb_n112, mult_msb_n111,
         mult_msb_n110, mult_msb_n109, mult_msb_n108, mult_msb_n107,
         mult_msb_n106, mult_msb_n105, mult_msb_n104, mult_msb_n103,
         mult_msb_n102, mult_msb_n101, mult_msb_n100, mult_msb_n99,
         mult_msb_n98, mult_msb_n97, mult_msb_n96, mult_msb_n95, mult_msb_n94,
         mult_msb_n93, mult_msb_n92, mult_msb_n91, mult_msb_n90, mult_msb_n89,
         mult_msb_n88, mult_msb_n87, mult_msb_n86, mult_msb_n85, mult_msb_n84,
         mult_msb_n83, mult_msb_n82, mult_msb_n81, mult_msb_n80, mult_msb_n79,
         mult_msb_n78, mult_msb_n77, mult_msb_n76, mult_msb_n75, mult_msb_n74,
         mult_msb_n73, mult_msb_n72, mult_msb_n71, mult_msb_n70, mult_msb_n69,
         mult_msb_n68, mult_msb_n67, mult_msb_n66, mult_msb_n65, mult_msb_n64,
         mult_msb_n63, mult_msb_n62, mult_msb_n61, mult_msb_n60, mult_msb_n59,
         mult_msb_n58, mult_msb_n57, mult_msb_n56, mult_msb_n55, mult_msb_n54,
         mult_msb_n53, mult_msb_n52, mult_msb_n51, mult_msb_n50, mult_msb_n49,
         mult_msb_n48, mult_msb_n47, mult_msb_n46, mult_msb_n45, mult_msb_n44,
         mult_msb_n43, mult_msb_n42, mult_msb_n41, mult_msb_n40, mult_msb_n39,
         mult_msb_n38, mult_msb_n37, mult_msb_n36, mult_msb_n35, mult_msb_n34,
         mult_msb_n33, mult_msb_Xi_mul_Yj_1__0_, mult_msb_Xi_mul_Yj_1__1_,
         mult_msb_Xi_mul_Yj_1__2_, mult_msb_Xi_mul_Yj_1__3_,
         mult_msb_Xi_mul_Yj_2__0_, mult_msb_Xi_mul_Yj_2__1_,
         mult_msb_Xi_mul_Yj_2__2_, mult_msb_Xi_mul_Yj_2__3_,
         mult_msb_Xi_mul_Yj_3__0_, mult_msb_Xi_mul_Yj_3__1_,
         mult_msb_Xi_mul_Yj_3__2_, mult_msb_Xi_mul_Yj_3__3_,
         mult_msb_Xi_mul_Yj_4__0_, mult_msb_Xi_mul_Yj_4__1_,
         mult_msb_Xi_mul_Yj_4__2_, mult_msb_Xi_mul_Yj_4__3_,
         mult_msb_Xi_mul_Yj_6__0_, mult_msb_Xi_mul_Yj_6__1_,
         mult_msb_Xi_mul_Yj_6__2_, mult_msb_Xi_mul_Yj_6__3_,
         mult_msb_Xi_mul_Yj_7__0_, mult_msb_Xi_mul_Yj_7__1_,
         mult_msb_Xi_mul_Yj_7__2_, mult_msb_Xi_mul_Yj_7__3_,
         mult_msb_Xi_mul_Yj_8__0_, mult_msb_Xi_mul_Yj_8__1_,
         mult_msb_Xi_mul_Yj_8__2_, mult_msb_Xi_mul_Yj_8__3_,
         mult_msb_Xi_mul_Yj_9__0_, mult_msb_Xi_mul_Yj_9__1_,
         mult_msb_Xi_mul_Yj_9__2_, mult_msb_Xi_mul_Yj_9__3_,
         mult_msb_Xi_mul_Yj_11__0_, mult_msb_Xi_mul_Yj_11__1_,
         mult_msb_Xi_mul_Yj_11__2_, mult_msb_Xi_mul_Yj_11__3_,
         mult_msb_Xi_mul_Yj_12__0_, mult_msb_Xi_mul_Yj_12__1_,
         mult_msb_Xi_mul_Yj_12__2_, mult_msb_Xi_mul_Yj_12__3_,
         mult_msb_Xi_mul_Yj_13__0_, mult_msb_Xi_mul_Yj_13__1_,
         mult_msb_Xi_mul_Yj_13__2_, mult_msb_Xi_mul_Yj_13__3_,
         mult_msb_Xi_mul_Yj_14__0_, mult_msb_Xi_mul_Yj_14__1_,
         mult_msb_Xi_mul_Yj_14__2_, mult_msb_Xi_mul_Yj_14__3_,
         mult_msb_gf4_mul_3_3_n77, mult_msb_gf4_mul_3_3_n76,
         mult_msb_gf4_mul_3_3_n75, mult_msb_gf4_mul_3_3_n74,
         mult_msb_gf4_mul_3_3_n73, mult_msb_gf4_mul_3_3_n72,
         mult_msb_gf4_mul_3_3_n71, mult_msb_gf4_mul_3_3_n70,
         mult_msb_gf4_mul_3_3_n69, mult_msb_gf4_mul_3_3_n68,
         mult_msb_gf4_mul_3_3_n67, mult_msb_gf4_mul_3_3_n66,
         mult_msb_gf4_mul_3_3_n65, mult_msb_gf4_mul_3_3_n64,
         mult_msb_gf4_mul_3_3_n63, mult_msb_gf4_mul_3_3_n62,
         mult_msb_gf4_mul_3_3_n61, mult_msb_gf4_mul_3_3_n60,
         mult_msb_gf4_mul_3_3_n59, mult_msb_gf4_mul_3_3_n58,
         mult_msb_gf4_mul_3_3_n57, mult_msb_gf4_mul_3_3_n56,
         mult_msb_gf4_mul_3_3_n55, mult_msb_gf4_mul_3_3_n54,
         mult_msb_gf4_mul_3_3_n53, mult_msb_gf4_mul_3_2_n77,
         mult_msb_gf4_mul_3_2_n76, mult_msb_gf4_mul_3_2_n75,
         mult_msb_gf4_mul_3_2_n74, mult_msb_gf4_mul_3_2_n73,
         mult_msb_gf4_mul_3_2_n72, mult_msb_gf4_mul_3_2_n71,
         mult_msb_gf4_mul_3_2_n70, mult_msb_gf4_mul_3_2_n69,
         mult_msb_gf4_mul_3_2_n68, mult_msb_gf4_mul_3_2_n67,
         mult_msb_gf4_mul_3_2_n66, mult_msb_gf4_mul_3_2_n65,
         mult_msb_gf4_mul_3_2_n64, mult_msb_gf4_mul_3_2_n63,
         mult_msb_gf4_mul_3_2_n62, mult_msb_gf4_mul_3_2_n61,
         mult_msb_gf4_mul_3_2_n60, mult_msb_gf4_mul_3_2_n59,
         mult_msb_gf4_mul_3_2_n58, mult_msb_gf4_mul_3_2_n57,
         mult_msb_gf4_mul_3_2_n56, mult_msb_gf4_mul_3_2_n55,
         mult_msb_gf4_mul_3_2_n54, mult_msb_gf4_mul_3_2_n53,
         mult_msb_gf4_mul_3_1_n77, mult_msb_gf4_mul_3_1_n76,
         mult_msb_gf4_mul_3_1_n75, mult_msb_gf4_mul_3_1_n74,
         mult_msb_gf4_mul_3_1_n73, mult_msb_gf4_mul_3_1_n72,
         mult_msb_gf4_mul_3_1_n71, mult_msb_gf4_mul_3_1_n70,
         mult_msb_gf4_mul_3_1_n69, mult_msb_gf4_mul_3_1_n68,
         mult_msb_gf4_mul_3_1_n67, mult_msb_gf4_mul_3_1_n66,
         mult_msb_gf4_mul_3_1_n65, mult_msb_gf4_mul_3_1_n64,
         mult_msb_gf4_mul_3_1_n63, mult_msb_gf4_mul_3_1_n62,
         mult_msb_gf4_mul_3_1_n61, mult_msb_gf4_mul_3_1_n60,
         mult_msb_gf4_mul_3_1_n59, mult_msb_gf4_mul_3_1_n58,
         mult_msb_gf4_mul_3_1_n57, mult_msb_gf4_mul_3_1_n56,
         mult_msb_gf4_mul_3_1_n55, mult_msb_gf4_mul_3_1_n54,
         mult_msb_gf4_mul_3_1_n53, mult_msb_gf4_mul_3_0_n77,
         mult_msb_gf4_mul_3_0_n76, mult_msb_gf4_mul_3_0_n75,
         mult_msb_gf4_mul_3_0_n74, mult_msb_gf4_mul_3_0_n73,
         mult_msb_gf4_mul_3_0_n72, mult_msb_gf4_mul_3_0_n71,
         mult_msb_gf4_mul_3_0_n70, mult_msb_gf4_mul_3_0_n69,
         mult_msb_gf4_mul_3_0_n68, mult_msb_gf4_mul_3_0_n67,
         mult_msb_gf4_mul_3_0_n66, mult_msb_gf4_mul_3_0_n65,
         mult_msb_gf4_mul_3_0_n64, mult_msb_gf4_mul_3_0_n63,
         mult_msb_gf4_mul_3_0_n62, mult_msb_gf4_mul_3_0_n61,
         mult_msb_gf4_mul_3_0_n60, mult_msb_gf4_mul_3_0_n59,
         mult_msb_gf4_mul_3_0_n58, mult_msb_gf4_mul_3_0_n57,
         mult_msb_gf4_mul_3_0_n56, mult_msb_gf4_mul_3_0_n55,
         mult_msb_gf4_mul_3_0_n54, mult_msb_gf4_mul_3_0_n53,
         mult_msb_gf4_mul_2_3_n77, mult_msb_gf4_mul_2_3_n76,
         mult_msb_gf4_mul_2_3_n75, mult_msb_gf4_mul_2_3_n74,
         mult_msb_gf4_mul_2_3_n73, mult_msb_gf4_mul_2_3_n72,
         mult_msb_gf4_mul_2_3_n71, mult_msb_gf4_mul_2_3_n70,
         mult_msb_gf4_mul_2_3_n69, mult_msb_gf4_mul_2_3_n68,
         mult_msb_gf4_mul_2_3_n67, mult_msb_gf4_mul_2_3_n66,
         mult_msb_gf4_mul_2_3_n65, mult_msb_gf4_mul_2_3_n64,
         mult_msb_gf4_mul_2_3_n63, mult_msb_gf4_mul_2_3_n62,
         mult_msb_gf4_mul_2_3_n61, mult_msb_gf4_mul_2_3_n60,
         mult_msb_gf4_mul_2_3_n59, mult_msb_gf4_mul_2_3_n58,
         mult_msb_gf4_mul_2_3_n57, mult_msb_gf4_mul_2_3_n56,
         mult_msb_gf4_mul_2_3_n55, mult_msb_gf4_mul_2_3_n54,
         mult_msb_gf4_mul_2_3_n53, mult_msb_gf4_mul_2_2_n77,
         mult_msb_gf4_mul_2_2_n76, mult_msb_gf4_mul_2_2_n75,
         mult_msb_gf4_mul_2_2_n74, mult_msb_gf4_mul_2_2_n73,
         mult_msb_gf4_mul_2_2_n72, mult_msb_gf4_mul_2_2_n71,
         mult_msb_gf4_mul_2_2_n70, mult_msb_gf4_mul_2_2_n69,
         mult_msb_gf4_mul_2_2_n68, mult_msb_gf4_mul_2_2_n67,
         mult_msb_gf4_mul_2_2_n66, mult_msb_gf4_mul_2_2_n65,
         mult_msb_gf4_mul_2_2_n64, mult_msb_gf4_mul_2_2_n63,
         mult_msb_gf4_mul_2_2_n62, mult_msb_gf4_mul_2_2_n61,
         mult_msb_gf4_mul_2_2_n60, mult_msb_gf4_mul_2_2_n59,
         mult_msb_gf4_mul_2_2_n58, mult_msb_gf4_mul_2_2_n57,
         mult_msb_gf4_mul_2_2_n56, mult_msb_gf4_mul_2_2_n55,
         mult_msb_gf4_mul_2_2_n54, mult_msb_gf4_mul_2_2_n53,
         mult_msb_gf4_mul_2_1_n77, mult_msb_gf4_mul_2_1_n76,
         mult_msb_gf4_mul_2_1_n75, mult_msb_gf4_mul_2_1_n74,
         mult_msb_gf4_mul_2_1_n73, mult_msb_gf4_mul_2_1_n72,
         mult_msb_gf4_mul_2_1_n71, mult_msb_gf4_mul_2_1_n70,
         mult_msb_gf4_mul_2_1_n69, mult_msb_gf4_mul_2_1_n68,
         mult_msb_gf4_mul_2_1_n67, mult_msb_gf4_mul_2_1_n66,
         mult_msb_gf4_mul_2_1_n65, mult_msb_gf4_mul_2_1_n64,
         mult_msb_gf4_mul_2_1_n63, mult_msb_gf4_mul_2_1_n62,
         mult_msb_gf4_mul_2_1_n61, mult_msb_gf4_mul_2_1_n60,
         mult_msb_gf4_mul_2_1_n59, mult_msb_gf4_mul_2_1_n58,
         mult_msb_gf4_mul_2_1_n57, mult_msb_gf4_mul_2_1_n56,
         mult_msb_gf4_mul_2_1_n55, mult_msb_gf4_mul_2_1_n54,
         mult_msb_gf4_mul_2_1_n53, mult_msb_gf4_mul_2_0_n77,
         mult_msb_gf4_mul_2_0_n76, mult_msb_gf4_mul_2_0_n75,
         mult_msb_gf4_mul_2_0_n74, mult_msb_gf4_mul_2_0_n73,
         mult_msb_gf4_mul_2_0_n72, mult_msb_gf4_mul_2_0_n71,
         mult_msb_gf4_mul_2_0_n70, mult_msb_gf4_mul_2_0_n69,
         mult_msb_gf4_mul_2_0_n68, mult_msb_gf4_mul_2_0_n67,
         mult_msb_gf4_mul_2_0_n66, mult_msb_gf4_mul_2_0_n65,
         mult_msb_gf4_mul_2_0_n64, mult_msb_gf4_mul_2_0_n63,
         mult_msb_gf4_mul_2_0_n62, mult_msb_gf4_mul_2_0_n61,
         mult_msb_gf4_mul_2_0_n60, mult_msb_gf4_mul_2_0_n59,
         mult_msb_gf4_mul_2_0_n58, mult_msb_gf4_mul_2_0_n57,
         mult_msb_gf4_mul_2_0_n56, mult_msb_gf4_mul_2_0_n55,
         mult_msb_gf4_mul_2_0_n54, mult_msb_gf4_mul_2_0_n53,
         mult_msb_gf4_mul_1_3_n77, mult_msb_gf4_mul_1_3_n76,
         mult_msb_gf4_mul_1_3_n75, mult_msb_gf4_mul_1_3_n74,
         mult_msb_gf4_mul_1_3_n73, mult_msb_gf4_mul_1_3_n72,
         mult_msb_gf4_mul_1_3_n71, mult_msb_gf4_mul_1_3_n70,
         mult_msb_gf4_mul_1_3_n69, mult_msb_gf4_mul_1_3_n68,
         mult_msb_gf4_mul_1_3_n67, mult_msb_gf4_mul_1_3_n66,
         mult_msb_gf4_mul_1_3_n65, mult_msb_gf4_mul_1_3_n64,
         mult_msb_gf4_mul_1_3_n63, mult_msb_gf4_mul_1_3_n62,
         mult_msb_gf4_mul_1_3_n61, mult_msb_gf4_mul_1_3_n60,
         mult_msb_gf4_mul_1_3_n59, mult_msb_gf4_mul_1_3_n58,
         mult_msb_gf4_mul_1_3_n57, mult_msb_gf4_mul_1_3_n56,
         mult_msb_gf4_mul_1_3_n55, mult_msb_gf4_mul_1_3_n54,
         mult_msb_gf4_mul_1_3_n53, mult_msb_gf4_mul_1_2_n77,
         mult_msb_gf4_mul_1_2_n76, mult_msb_gf4_mul_1_2_n75,
         mult_msb_gf4_mul_1_2_n74, mult_msb_gf4_mul_1_2_n73,
         mult_msb_gf4_mul_1_2_n72, mult_msb_gf4_mul_1_2_n71,
         mult_msb_gf4_mul_1_2_n70, mult_msb_gf4_mul_1_2_n69,
         mult_msb_gf4_mul_1_2_n68, mult_msb_gf4_mul_1_2_n67,
         mult_msb_gf4_mul_1_2_n66, mult_msb_gf4_mul_1_2_n65,
         mult_msb_gf4_mul_1_2_n64, mult_msb_gf4_mul_1_2_n63,
         mult_msb_gf4_mul_1_2_n62, mult_msb_gf4_mul_1_2_n61,
         mult_msb_gf4_mul_1_2_n60, mult_msb_gf4_mul_1_2_n59,
         mult_msb_gf4_mul_1_2_n58, mult_msb_gf4_mul_1_2_n57,
         mult_msb_gf4_mul_1_2_n56, mult_msb_gf4_mul_1_2_n55,
         mult_msb_gf4_mul_1_2_n54, mult_msb_gf4_mul_1_2_n53,
         mult_msb_gf4_mul_1_1_n77, mult_msb_gf4_mul_1_1_n76,
         mult_msb_gf4_mul_1_1_n75, mult_msb_gf4_mul_1_1_n74,
         mult_msb_gf4_mul_1_1_n73, mult_msb_gf4_mul_1_1_n72,
         mult_msb_gf4_mul_1_1_n71, mult_msb_gf4_mul_1_1_n70,
         mult_msb_gf4_mul_1_1_n69, mult_msb_gf4_mul_1_1_n68,
         mult_msb_gf4_mul_1_1_n67, mult_msb_gf4_mul_1_1_n66,
         mult_msb_gf4_mul_1_1_n65, mult_msb_gf4_mul_1_1_n64,
         mult_msb_gf4_mul_1_1_n63, mult_msb_gf4_mul_1_1_n62,
         mult_msb_gf4_mul_1_1_n61, mult_msb_gf4_mul_1_1_n60,
         mult_msb_gf4_mul_1_1_n59, mult_msb_gf4_mul_1_1_n58,
         mult_msb_gf4_mul_1_1_n57, mult_msb_gf4_mul_1_1_n56,
         mult_msb_gf4_mul_1_1_n55, mult_msb_gf4_mul_1_1_n54,
         mult_msb_gf4_mul_1_1_n53, mult_msb_gf4_mul_1_0_n77,
         mult_msb_gf4_mul_1_0_n76, mult_msb_gf4_mul_1_0_n75,
         mult_msb_gf4_mul_1_0_n74, mult_msb_gf4_mul_1_0_n73,
         mult_msb_gf4_mul_1_0_n72, mult_msb_gf4_mul_1_0_n71,
         mult_msb_gf4_mul_1_0_n70, mult_msb_gf4_mul_1_0_n69,
         mult_msb_gf4_mul_1_0_n68, mult_msb_gf4_mul_1_0_n67,
         mult_msb_gf4_mul_1_0_n66, mult_msb_gf4_mul_1_0_n65,
         mult_msb_gf4_mul_1_0_n64, mult_msb_gf4_mul_1_0_n63,
         mult_msb_gf4_mul_1_0_n62, mult_msb_gf4_mul_1_0_n61,
         mult_msb_gf4_mul_1_0_n60, mult_msb_gf4_mul_1_0_n59,
         mult_msb_gf4_mul_1_0_n58, mult_msb_gf4_mul_1_0_n57,
         mult_msb_gf4_mul_1_0_n56, mult_msb_gf4_mul_1_0_n55,
         mult_msb_gf4_mul_1_0_n54, mult_msb_gf4_mul_1_0_n53,
         mult_msb_gf4_mul_0_3_n77, mult_msb_gf4_mul_0_3_n76,
         mult_msb_gf4_mul_0_3_n75, mult_msb_gf4_mul_0_3_n74,
         mult_msb_gf4_mul_0_3_n73, mult_msb_gf4_mul_0_3_n72,
         mult_msb_gf4_mul_0_3_n71, mult_msb_gf4_mul_0_3_n70,
         mult_msb_gf4_mul_0_3_n69, mult_msb_gf4_mul_0_3_n68,
         mult_msb_gf4_mul_0_3_n67, mult_msb_gf4_mul_0_3_n66,
         mult_msb_gf4_mul_0_3_n65, mult_msb_gf4_mul_0_3_n64,
         mult_msb_gf4_mul_0_3_n63, mult_msb_gf4_mul_0_3_n62,
         mult_msb_gf4_mul_0_3_n61, mult_msb_gf4_mul_0_3_n60,
         mult_msb_gf4_mul_0_3_n59, mult_msb_gf4_mul_0_3_n58,
         mult_msb_gf4_mul_0_3_n57, mult_msb_gf4_mul_0_3_n56,
         mult_msb_gf4_mul_0_3_n55, mult_msb_gf4_mul_0_3_n54,
         mult_msb_gf4_mul_0_3_n53, mult_msb_gf4_mul_0_2_n77,
         mult_msb_gf4_mul_0_2_n76, mult_msb_gf4_mul_0_2_n75,
         mult_msb_gf4_mul_0_2_n74, mult_msb_gf4_mul_0_2_n73,
         mult_msb_gf4_mul_0_2_n72, mult_msb_gf4_mul_0_2_n71,
         mult_msb_gf4_mul_0_2_n70, mult_msb_gf4_mul_0_2_n69,
         mult_msb_gf4_mul_0_2_n68, mult_msb_gf4_mul_0_2_n67,
         mult_msb_gf4_mul_0_2_n66, mult_msb_gf4_mul_0_2_n65,
         mult_msb_gf4_mul_0_2_n64, mult_msb_gf4_mul_0_2_n63,
         mult_msb_gf4_mul_0_2_n62, mult_msb_gf4_mul_0_2_n61,
         mult_msb_gf4_mul_0_2_n60, mult_msb_gf4_mul_0_2_n59,
         mult_msb_gf4_mul_0_2_n58, mult_msb_gf4_mul_0_2_n57,
         mult_msb_gf4_mul_0_2_n56, mult_msb_gf4_mul_0_2_n55,
         mult_msb_gf4_mul_0_2_n54, mult_msb_gf4_mul_0_2_n53,
         mult_msb_gf4_mul_0_1_n77, mult_msb_gf4_mul_0_1_n76,
         mult_msb_gf4_mul_0_1_n75, mult_msb_gf4_mul_0_1_n74,
         mult_msb_gf4_mul_0_1_n73, mult_msb_gf4_mul_0_1_n72,
         mult_msb_gf4_mul_0_1_n71, mult_msb_gf4_mul_0_1_n70,
         mult_msb_gf4_mul_0_1_n69, mult_msb_gf4_mul_0_1_n68,
         mult_msb_gf4_mul_0_1_n67, mult_msb_gf4_mul_0_1_n66,
         mult_msb_gf4_mul_0_1_n65, mult_msb_gf4_mul_0_1_n64,
         mult_msb_gf4_mul_0_1_n63, mult_msb_gf4_mul_0_1_n62,
         mult_msb_gf4_mul_0_1_n61, mult_msb_gf4_mul_0_1_n60,
         mult_msb_gf4_mul_0_1_n59, mult_msb_gf4_mul_0_1_n58,
         mult_msb_gf4_mul_0_1_n57, mult_msb_gf4_mul_0_1_n56,
         mult_msb_gf4_mul_0_1_n55, mult_msb_gf4_mul_0_1_n54,
         mult_msb_gf4_mul_0_1_n53, mult_msb_gf4_mul_0_0_n77,
         mult_msb_gf4_mul_0_0_n76, mult_msb_gf4_mul_0_0_n75,
         mult_msb_gf4_mul_0_0_n74, mult_msb_gf4_mul_0_0_n73,
         mult_msb_gf4_mul_0_0_n72, mult_msb_gf4_mul_0_0_n71,
         mult_msb_gf4_mul_0_0_n70, mult_msb_gf4_mul_0_0_n69,
         mult_msb_gf4_mul_0_0_n68, mult_msb_gf4_mul_0_0_n67,
         mult_msb_gf4_mul_0_0_n66, mult_msb_gf4_mul_0_0_n65,
         mult_msb_gf4_mul_0_0_n64, mult_msb_gf4_mul_0_0_n63,
         mult_msb_gf4_mul_0_0_n62, mult_msb_gf4_mul_0_0_n61,
         mult_msb_gf4_mul_0_0_n60, mult_msb_gf4_mul_0_0_n59,
         mult_msb_gf4_mul_0_0_n58, mult_msb_gf4_mul_0_0_n57,
         mult_msb_gf4_mul_0_0_n56, mult_msb_gf4_mul_0_0_n55,
         mult_msb_gf4_mul_0_0_n54, mult_msb_gf4_mul_0_0_n53, mult_lsb_n128,
         mult_lsb_n127, mult_lsb_n126, mult_lsb_n125, mult_lsb_n124,
         mult_lsb_n123, mult_lsb_n122, mult_lsb_n121, mult_lsb_n120,
         mult_lsb_n119, mult_lsb_n118, mult_lsb_n117, mult_lsb_n116,
         mult_lsb_n115, mult_lsb_n114, mult_lsb_n113, mult_lsb_n112,
         mult_lsb_n111, mult_lsb_n110, mult_lsb_n109, mult_lsb_n108,
         mult_lsb_n107, mult_lsb_n106, mult_lsb_n105, mult_lsb_n104,
         mult_lsb_n103, mult_lsb_n102, mult_lsb_n101, mult_lsb_n100,
         mult_lsb_n99, mult_lsb_n98, mult_lsb_n97, mult_lsb_n96, mult_lsb_n95,
         mult_lsb_n94, mult_lsb_n93, mult_lsb_n92, mult_lsb_n91, mult_lsb_n90,
         mult_lsb_n89, mult_lsb_n88, mult_lsb_n87, mult_lsb_n86, mult_lsb_n85,
         mult_lsb_n84, mult_lsb_n83, mult_lsb_n82, mult_lsb_n81, mult_lsb_n80,
         mult_lsb_n79, mult_lsb_n78, mult_lsb_n77, mult_lsb_n76, mult_lsb_n75,
         mult_lsb_n74, mult_lsb_n73, mult_lsb_n72, mult_lsb_n71, mult_lsb_n70,
         mult_lsb_n69, mult_lsb_n68, mult_lsb_n67, mult_lsb_n66, mult_lsb_n65,
         mult_lsb_n64, mult_lsb_n63, mult_lsb_n62, mult_lsb_n61, mult_lsb_n60,
         mult_lsb_n59, mult_lsb_n58, mult_lsb_n57, mult_lsb_n56, mult_lsb_n55,
         mult_lsb_n54, mult_lsb_n53, mult_lsb_n52, mult_lsb_n51, mult_lsb_n50,
         mult_lsb_n49, mult_lsb_n48, mult_lsb_n47, mult_lsb_n46, mult_lsb_n45,
         mult_lsb_n44, mult_lsb_n43, mult_lsb_n42, mult_lsb_n41, mult_lsb_n40,
         mult_lsb_n39, mult_lsb_n38, mult_lsb_n37, mult_lsb_n36, mult_lsb_n35,
         mult_lsb_n34, mult_lsb_n33, mult_lsb_Xi_mul_Yj_1__0_,
         mult_lsb_Xi_mul_Yj_1__1_, mult_lsb_Xi_mul_Yj_1__2_,
         mult_lsb_Xi_mul_Yj_1__3_, mult_lsb_Xi_mul_Yj_2__0_,
         mult_lsb_Xi_mul_Yj_2__1_, mult_lsb_Xi_mul_Yj_2__2_,
         mult_lsb_Xi_mul_Yj_2__3_, mult_lsb_Xi_mul_Yj_3__0_,
         mult_lsb_Xi_mul_Yj_3__1_, mult_lsb_Xi_mul_Yj_3__2_,
         mult_lsb_Xi_mul_Yj_3__3_, mult_lsb_Xi_mul_Yj_4__0_,
         mult_lsb_Xi_mul_Yj_4__1_, mult_lsb_Xi_mul_Yj_4__2_,
         mult_lsb_Xi_mul_Yj_4__3_, mult_lsb_Xi_mul_Yj_6__0_,
         mult_lsb_Xi_mul_Yj_6__1_, mult_lsb_Xi_mul_Yj_6__2_,
         mult_lsb_Xi_mul_Yj_6__3_, mult_lsb_Xi_mul_Yj_7__0_,
         mult_lsb_Xi_mul_Yj_7__1_, mult_lsb_Xi_mul_Yj_7__2_,
         mult_lsb_Xi_mul_Yj_7__3_, mult_lsb_Xi_mul_Yj_8__0_,
         mult_lsb_Xi_mul_Yj_8__1_, mult_lsb_Xi_mul_Yj_8__2_,
         mult_lsb_Xi_mul_Yj_8__3_, mult_lsb_Xi_mul_Yj_9__0_,
         mult_lsb_Xi_mul_Yj_9__1_, mult_lsb_Xi_mul_Yj_9__2_,
         mult_lsb_Xi_mul_Yj_9__3_, mult_lsb_Xi_mul_Yj_11__0_,
         mult_lsb_Xi_mul_Yj_11__1_, mult_lsb_Xi_mul_Yj_11__2_,
         mult_lsb_Xi_mul_Yj_11__3_, mult_lsb_Xi_mul_Yj_12__0_,
         mult_lsb_Xi_mul_Yj_12__1_, mult_lsb_Xi_mul_Yj_12__2_,
         mult_lsb_Xi_mul_Yj_12__3_, mult_lsb_Xi_mul_Yj_13__0_,
         mult_lsb_Xi_mul_Yj_13__1_, mult_lsb_Xi_mul_Yj_13__2_,
         mult_lsb_Xi_mul_Yj_13__3_, mult_lsb_Xi_mul_Yj_14__0_,
         mult_lsb_Xi_mul_Yj_14__1_, mult_lsb_Xi_mul_Yj_14__2_,
         mult_lsb_Xi_mul_Yj_14__3_, mult_lsb_gf4_mul_3_3_n77,
         mult_lsb_gf4_mul_3_3_n76, mult_lsb_gf4_mul_3_3_n75,
         mult_lsb_gf4_mul_3_3_n74, mult_lsb_gf4_mul_3_3_n73,
         mult_lsb_gf4_mul_3_3_n72, mult_lsb_gf4_mul_3_3_n71,
         mult_lsb_gf4_mul_3_3_n70, mult_lsb_gf4_mul_3_3_n69,
         mult_lsb_gf4_mul_3_3_n68, mult_lsb_gf4_mul_3_3_n67,
         mult_lsb_gf4_mul_3_3_n66, mult_lsb_gf4_mul_3_3_n65,
         mult_lsb_gf4_mul_3_3_n64, mult_lsb_gf4_mul_3_3_n63,
         mult_lsb_gf4_mul_3_3_n62, mult_lsb_gf4_mul_3_3_n61,
         mult_lsb_gf4_mul_3_3_n60, mult_lsb_gf4_mul_3_3_n59,
         mult_lsb_gf4_mul_3_3_n58, mult_lsb_gf4_mul_3_3_n57,
         mult_lsb_gf4_mul_3_3_n56, mult_lsb_gf4_mul_3_3_n55,
         mult_lsb_gf4_mul_3_3_n54, mult_lsb_gf4_mul_3_3_n53,
         mult_lsb_gf4_mul_3_2_n77, mult_lsb_gf4_mul_3_2_n76,
         mult_lsb_gf4_mul_3_2_n75, mult_lsb_gf4_mul_3_2_n74,
         mult_lsb_gf4_mul_3_2_n73, mult_lsb_gf4_mul_3_2_n72,
         mult_lsb_gf4_mul_3_2_n71, mult_lsb_gf4_mul_3_2_n70,
         mult_lsb_gf4_mul_3_2_n69, mult_lsb_gf4_mul_3_2_n68,
         mult_lsb_gf4_mul_3_2_n67, mult_lsb_gf4_mul_3_2_n66,
         mult_lsb_gf4_mul_3_2_n65, mult_lsb_gf4_mul_3_2_n64,
         mult_lsb_gf4_mul_3_2_n63, mult_lsb_gf4_mul_3_2_n62,
         mult_lsb_gf4_mul_3_2_n61, mult_lsb_gf4_mul_3_2_n60,
         mult_lsb_gf4_mul_3_2_n59, mult_lsb_gf4_mul_3_2_n58,
         mult_lsb_gf4_mul_3_2_n57, mult_lsb_gf4_mul_3_2_n56,
         mult_lsb_gf4_mul_3_2_n55, mult_lsb_gf4_mul_3_2_n54,
         mult_lsb_gf4_mul_3_2_n53, mult_lsb_gf4_mul_3_1_n77,
         mult_lsb_gf4_mul_3_1_n76, mult_lsb_gf4_mul_3_1_n75,
         mult_lsb_gf4_mul_3_1_n74, mult_lsb_gf4_mul_3_1_n73,
         mult_lsb_gf4_mul_3_1_n72, mult_lsb_gf4_mul_3_1_n71,
         mult_lsb_gf4_mul_3_1_n70, mult_lsb_gf4_mul_3_1_n69,
         mult_lsb_gf4_mul_3_1_n68, mult_lsb_gf4_mul_3_1_n67,
         mult_lsb_gf4_mul_3_1_n66, mult_lsb_gf4_mul_3_1_n65,
         mult_lsb_gf4_mul_3_1_n64, mult_lsb_gf4_mul_3_1_n63,
         mult_lsb_gf4_mul_3_1_n62, mult_lsb_gf4_mul_3_1_n61,
         mult_lsb_gf4_mul_3_1_n60, mult_lsb_gf4_mul_3_1_n59,
         mult_lsb_gf4_mul_3_1_n58, mult_lsb_gf4_mul_3_1_n57,
         mult_lsb_gf4_mul_3_1_n56, mult_lsb_gf4_mul_3_1_n55,
         mult_lsb_gf4_mul_3_1_n54, mult_lsb_gf4_mul_3_1_n53,
         mult_lsb_gf4_mul_3_0_n77, mult_lsb_gf4_mul_3_0_n76,
         mult_lsb_gf4_mul_3_0_n75, mult_lsb_gf4_mul_3_0_n74,
         mult_lsb_gf4_mul_3_0_n73, mult_lsb_gf4_mul_3_0_n72,
         mult_lsb_gf4_mul_3_0_n71, mult_lsb_gf4_mul_3_0_n70,
         mult_lsb_gf4_mul_3_0_n69, mult_lsb_gf4_mul_3_0_n68,
         mult_lsb_gf4_mul_3_0_n67, mult_lsb_gf4_mul_3_0_n66,
         mult_lsb_gf4_mul_3_0_n65, mult_lsb_gf4_mul_3_0_n64,
         mult_lsb_gf4_mul_3_0_n63, mult_lsb_gf4_mul_3_0_n62,
         mult_lsb_gf4_mul_3_0_n61, mult_lsb_gf4_mul_3_0_n60,
         mult_lsb_gf4_mul_3_0_n59, mult_lsb_gf4_mul_3_0_n58,
         mult_lsb_gf4_mul_3_0_n57, mult_lsb_gf4_mul_3_0_n56,
         mult_lsb_gf4_mul_3_0_n55, mult_lsb_gf4_mul_3_0_n54,
         mult_lsb_gf4_mul_3_0_n53, mult_lsb_gf4_mul_2_3_n77,
         mult_lsb_gf4_mul_2_3_n76, mult_lsb_gf4_mul_2_3_n75,
         mult_lsb_gf4_mul_2_3_n74, mult_lsb_gf4_mul_2_3_n73,
         mult_lsb_gf4_mul_2_3_n72, mult_lsb_gf4_mul_2_3_n71,
         mult_lsb_gf4_mul_2_3_n70, mult_lsb_gf4_mul_2_3_n69,
         mult_lsb_gf4_mul_2_3_n68, mult_lsb_gf4_mul_2_3_n67,
         mult_lsb_gf4_mul_2_3_n66, mult_lsb_gf4_mul_2_3_n65,
         mult_lsb_gf4_mul_2_3_n64, mult_lsb_gf4_mul_2_3_n63,
         mult_lsb_gf4_mul_2_3_n62, mult_lsb_gf4_mul_2_3_n61,
         mult_lsb_gf4_mul_2_3_n60, mult_lsb_gf4_mul_2_3_n59,
         mult_lsb_gf4_mul_2_3_n58, mult_lsb_gf4_mul_2_3_n57,
         mult_lsb_gf4_mul_2_3_n56, mult_lsb_gf4_mul_2_3_n55,
         mult_lsb_gf4_mul_2_3_n54, mult_lsb_gf4_mul_2_3_n53,
         mult_lsb_gf4_mul_2_2_n77, mult_lsb_gf4_mul_2_2_n76,
         mult_lsb_gf4_mul_2_2_n75, mult_lsb_gf4_mul_2_2_n74,
         mult_lsb_gf4_mul_2_2_n73, mult_lsb_gf4_mul_2_2_n72,
         mult_lsb_gf4_mul_2_2_n71, mult_lsb_gf4_mul_2_2_n70,
         mult_lsb_gf4_mul_2_2_n69, mult_lsb_gf4_mul_2_2_n68,
         mult_lsb_gf4_mul_2_2_n67, mult_lsb_gf4_mul_2_2_n66,
         mult_lsb_gf4_mul_2_2_n65, mult_lsb_gf4_mul_2_2_n64,
         mult_lsb_gf4_mul_2_2_n63, mult_lsb_gf4_mul_2_2_n62,
         mult_lsb_gf4_mul_2_2_n61, mult_lsb_gf4_mul_2_2_n60,
         mult_lsb_gf4_mul_2_2_n59, mult_lsb_gf4_mul_2_2_n58,
         mult_lsb_gf4_mul_2_2_n57, mult_lsb_gf4_mul_2_2_n56,
         mult_lsb_gf4_mul_2_2_n55, mult_lsb_gf4_mul_2_2_n54,
         mult_lsb_gf4_mul_2_2_n53, mult_lsb_gf4_mul_2_1_n77,
         mult_lsb_gf4_mul_2_1_n76, mult_lsb_gf4_mul_2_1_n75,
         mult_lsb_gf4_mul_2_1_n74, mult_lsb_gf4_mul_2_1_n73,
         mult_lsb_gf4_mul_2_1_n72, mult_lsb_gf4_mul_2_1_n71,
         mult_lsb_gf4_mul_2_1_n70, mult_lsb_gf4_mul_2_1_n69,
         mult_lsb_gf4_mul_2_1_n68, mult_lsb_gf4_mul_2_1_n67,
         mult_lsb_gf4_mul_2_1_n66, mult_lsb_gf4_mul_2_1_n65,
         mult_lsb_gf4_mul_2_1_n64, mult_lsb_gf4_mul_2_1_n63,
         mult_lsb_gf4_mul_2_1_n62, mult_lsb_gf4_mul_2_1_n61,
         mult_lsb_gf4_mul_2_1_n60, mult_lsb_gf4_mul_2_1_n59,
         mult_lsb_gf4_mul_2_1_n58, mult_lsb_gf4_mul_2_1_n57,
         mult_lsb_gf4_mul_2_1_n56, mult_lsb_gf4_mul_2_1_n55,
         mult_lsb_gf4_mul_2_1_n54, mult_lsb_gf4_mul_2_1_n53,
         mult_lsb_gf4_mul_2_0_n77, mult_lsb_gf4_mul_2_0_n76,
         mult_lsb_gf4_mul_2_0_n75, mult_lsb_gf4_mul_2_0_n74,
         mult_lsb_gf4_mul_2_0_n73, mult_lsb_gf4_mul_2_0_n72,
         mult_lsb_gf4_mul_2_0_n71, mult_lsb_gf4_mul_2_0_n70,
         mult_lsb_gf4_mul_2_0_n69, mult_lsb_gf4_mul_2_0_n68,
         mult_lsb_gf4_mul_2_0_n67, mult_lsb_gf4_mul_2_0_n66,
         mult_lsb_gf4_mul_2_0_n65, mult_lsb_gf4_mul_2_0_n64,
         mult_lsb_gf4_mul_2_0_n63, mult_lsb_gf4_mul_2_0_n62,
         mult_lsb_gf4_mul_2_0_n61, mult_lsb_gf4_mul_2_0_n60,
         mult_lsb_gf4_mul_2_0_n59, mult_lsb_gf4_mul_2_0_n58,
         mult_lsb_gf4_mul_2_0_n57, mult_lsb_gf4_mul_2_0_n56,
         mult_lsb_gf4_mul_2_0_n55, mult_lsb_gf4_mul_2_0_n54,
         mult_lsb_gf4_mul_2_0_n53, mult_lsb_gf4_mul_1_3_n77,
         mult_lsb_gf4_mul_1_3_n76, mult_lsb_gf4_mul_1_3_n75,
         mult_lsb_gf4_mul_1_3_n74, mult_lsb_gf4_mul_1_3_n73,
         mult_lsb_gf4_mul_1_3_n72, mult_lsb_gf4_mul_1_3_n71,
         mult_lsb_gf4_mul_1_3_n70, mult_lsb_gf4_mul_1_3_n69,
         mult_lsb_gf4_mul_1_3_n68, mult_lsb_gf4_mul_1_3_n67,
         mult_lsb_gf4_mul_1_3_n66, mult_lsb_gf4_mul_1_3_n65,
         mult_lsb_gf4_mul_1_3_n64, mult_lsb_gf4_mul_1_3_n63,
         mult_lsb_gf4_mul_1_3_n62, mult_lsb_gf4_mul_1_3_n61,
         mult_lsb_gf4_mul_1_3_n60, mult_lsb_gf4_mul_1_3_n59,
         mult_lsb_gf4_mul_1_3_n58, mult_lsb_gf4_mul_1_3_n57,
         mult_lsb_gf4_mul_1_3_n56, mult_lsb_gf4_mul_1_3_n55,
         mult_lsb_gf4_mul_1_3_n54, mult_lsb_gf4_mul_1_3_n53,
         mult_lsb_gf4_mul_1_2_n77, mult_lsb_gf4_mul_1_2_n76,
         mult_lsb_gf4_mul_1_2_n75, mult_lsb_gf4_mul_1_2_n74,
         mult_lsb_gf4_mul_1_2_n73, mult_lsb_gf4_mul_1_2_n72,
         mult_lsb_gf4_mul_1_2_n71, mult_lsb_gf4_mul_1_2_n70,
         mult_lsb_gf4_mul_1_2_n69, mult_lsb_gf4_mul_1_2_n68,
         mult_lsb_gf4_mul_1_2_n67, mult_lsb_gf4_mul_1_2_n66,
         mult_lsb_gf4_mul_1_2_n65, mult_lsb_gf4_mul_1_2_n64,
         mult_lsb_gf4_mul_1_2_n63, mult_lsb_gf4_mul_1_2_n62,
         mult_lsb_gf4_mul_1_2_n61, mult_lsb_gf4_mul_1_2_n60,
         mult_lsb_gf4_mul_1_2_n59, mult_lsb_gf4_mul_1_2_n58,
         mult_lsb_gf4_mul_1_2_n57, mult_lsb_gf4_mul_1_2_n56,
         mult_lsb_gf4_mul_1_2_n55, mult_lsb_gf4_mul_1_2_n54,
         mult_lsb_gf4_mul_1_2_n53, mult_lsb_gf4_mul_1_1_n77,
         mult_lsb_gf4_mul_1_1_n76, mult_lsb_gf4_mul_1_1_n75,
         mult_lsb_gf4_mul_1_1_n74, mult_lsb_gf4_mul_1_1_n73,
         mult_lsb_gf4_mul_1_1_n72, mult_lsb_gf4_mul_1_1_n71,
         mult_lsb_gf4_mul_1_1_n70, mult_lsb_gf4_mul_1_1_n69,
         mult_lsb_gf4_mul_1_1_n68, mult_lsb_gf4_mul_1_1_n67,
         mult_lsb_gf4_mul_1_1_n66, mult_lsb_gf4_mul_1_1_n65,
         mult_lsb_gf4_mul_1_1_n64, mult_lsb_gf4_mul_1_1_n63,
         mult_lsb_gf4_mul_1_1_n62, mult_lsb_gf4_mul_1_1_n61,
         mult_lsb_gf4_mul_1_1_n60, mult_lsb_gf4_mul_1_1_n59,
         mult_lsb_gf4_mul_1_1_n58, mult_lsb_gf4_mul_1_1_n57,
         mult_lsb_gf4_mul_1_1_n56, mult_lsb_gf4_mul_1_1_n55,
         mult_lsb_gf4_mul_1_1_n54, mult_lsb_gf4_mul_1_1_n53,
         mult_lsb_gf4_mul_1_0_n77, mult_lsb_gf4_mul_1_0_n76,
         mult_lsb_gf4_mul_1_0_n75, mult_lsb_gf4_mul_1_0_n74,
         mult_lsb_gf4_mul_1_0_n73, mult_lsb_gf4_mul_1_0_n72,
         mult_lsb_gf4_mul_1_0_n71, mult_lsb_gf4_mul_1_0_n70,
         mult_lsb_gf4_mul_1_0_n69, mult_lsb_gf4_mul_1_0_n68,
         mult_lsb_gf4_mul_1_0_n67, mult_lsb_gf4_mul_1_0_n66,
         mult_lsb_gf4_mul_1_0_n65, mult_lsb_gf4_mul_1_0_n64,
         mult_lsb_gf4_mul_1_0_n63, mult_lsb_gf4_mul_1_0_n62,
         mult_lsb_gf4_mul_1_0_n61, mult_lsb_gf4_mul_1_0_n60,
         mult_lsb_gf4_mul_1_0_n59, mult_lsb_gf4_mul_1_0_n58,
         mult_lsb_gf4_mul_1_0_n57, mult_lsb_gf4_mul_1_0_n56,
         mult_lsb_gf4_mul_1_0_n55, mult_lsb_gf4_mul_1_0_n54,
         mult_lsb_gf4_mul_1_0_n53, mult_lsb_gf4_mul_0_3_n77,
         mult_lsb_gf4_mul_0_3_n76, mult_lsb_gf4_mul_0_3_n75,
         mult_lsb_gf4_mul_0_3_n74, mult_lsb_gf4_mul_0_3_n73,
         mult_lsb_gf4_mul_0_3_n72, mult_lsb_gf4_mul_0_3_n71,
         mult_lsb_gf4_mul_0_3_n70, mult_lsb_gf4_mul_0_3_n69,
         mult_lsb_gf4_mul_0_3_n68, mult_lsb_gf4_mul_0_3_n67,
         mult_lsb_gf4_mul_0_3_n66, mult_lsb_gf4_mul_0_3_n65,
         mult_lsb_gf4_mul_0_3_n64, mult_lsb_gf4_mul_0_3_n63,
         mult_lsb_gf4_mul_0_3_n62, mult_lsb_gf4_mul_0_3_n61,
         mult_lsb_gf4_mul_0_3_n60, mult_lsb_gf4_mul_0_3_n59,
         mult_lsb_gf4_mul_0_3_n58, mult_lsb_gf4_mul_0_3_n57,
         mult_lsb_gf4_mul_0_3_n56, mult_lsb_gf4_mul_0_3_n55,
         mult_lsb_gf4_mul_0_3_n54, mult_lsb_gf4_mul_0_3_n53,
         mult_lsb_gf4_mul_0_2_n77, mult_lsb_gf4_mul_0_2_n76,
         mult_lsb_gf4_mul_0_2_n75, mult_lsb_gf4_mul_0_2_n74,
         mult_lsb_gf4_mul_0_2_n73, mult_lsb_gf4_mul_0_2_n72,
         mult_lsb_gf4_mul_0_2_n71, mult_lsb_gf4_mul_0_2_n70,
         mult_lsb_gf4_mul_0_2_n69, mult_lsb_gf4_mul_0_2_n68,
         mult_lsb_gf4_mul_0_2_n67, mult_lsb_gf4_mul_0_2_n66,
         mult_lsb_gf4_mul_0_2_n65, mult_lsb_gf4_mul_0_2_n64,
         mult_lsb_gf4_mul_0_2_n63, mult_lsb_gf4_mul_0_2_n62,
         mult_lsb_gf4_mul_0_2_n61, mult_lsb_gf4_mul_0_2_n60,
         mult_lsb_gf4_mul_0_2_n59, mult_lsb_gf4_mul_0_2_n58,
         mult_lsb_gf4_mul_0_2_n57, mult_lsb_gf4_mul_0_2_n56,
         mult_lsb_gf4_mul_0_2_n55, mult_lsb_gf4_mul_0_2_n54,
         mult_lsb_gf4_mul_0_2_n53, mult_lsb_gf4_mul_0_1_n77,
         mult_lsb_gf4_mul_0_1_n76, mult_lsb_gf4_mul_0_1_n75,
         mult_lsb_gf4_mul_0_1_n74, mult_lsb_gf4_mul_0_1_n73,
         mult_lsb_gf4_mul_0_1_n72, mult_lsb_gf4_mul_0_1_n71,
         mult_lsb_gf4_mul_0_1_n70, mult_lsb_gf4_mul_0_1_n69,
         mult_lsb_gf4_mul_0_1_n68, mult_lsb_gf4_mul_0_1_n67,
         mult_lsb_gf4_mul_0_1_n66, mult_lsb_gf4_mul_0_1_n65,
         mult_lsb_gf4_mul_0_1_n64, mult_lsb_gf4_mul_0_1_n63,
         mult_lsb_gf4_mul_0_1_n62, mult_lsb_gf4_mul_0_1_n61,
         mult_lsb_gf4_mul_0_1_n60, mult_lsb_gf4_mul_0_1_n59,
         mult_lsb_gf4_mul_0_1_n58, mult_lsb_gf4_mul_0_1_n57,
         mult_lsb_gf4_mul_0_1_n56, mult_lsb_gf4_mul_0_1_n55,
         mult_lsb_gf4_mul_0_1_n54, mult_lsb_gf4_mul_0_1_n53,
         mult_lsb_gf4_mul_0_0_n77, mult_lsb_gf4_mul_0_0_n76,
         mult_lsb_gf4_mul_0_0_n75, mult_lsb_gf4_mul_0_0_n74,
         mult_lsb_gf4_mul_0_0_n73, mult_lsb_gf4_mul_0_0_n72,
         mult_lsb_gf4_mul_0_0_n71, mult_lsb_gf4_mul_0_0_n70,
         mult_lsb_gf4_mul_0_0_n69, mult_lsb_gf4_mul_0_0_n68,
         mult_lsb_gf4_mul_0_0_n67, mult_lsb_gf4_mul_0_0_n66,
         mult_lsb_gf4_mul_0_0_n65, mult_lsb_gf4_mul_0_0_n64,
         mult_lsb_gf4_mul_0_0_n63, mult_lsb_gf4_mul_0_0_n62,
         mult_lsb_gf4_mul_0_0_n61, mult_lsb_gf4_mul_0_0_n60,
         mult_lsb_gf4_mul_0_0_n59, mult_lsb_gf4_mul_0_0_n58,
         mult_lsb_gf4_mul_0_0_n57, mult_lsb_gf4_mul_0_0_n56,
         mult_lsb_gf4_mul_0_0_n55, mult_lsb_gf4_mul_0_0_n54,
         mult_lsb_gf4_mul_0_0_n53;
  wire   [15:0] Y1xD;
  wire   [15:0] Y0xD;
  wire   [15:0] InverterInxDP;
  wire   [15:0] InverterInxD;
  wire   [15:0] Y0_0xDP;
  wire   [15:0] Y0_1xDP;
  wire   [15:0] Y0_2xDP;
  wire   [15:0] Y0_3xDP;
  wire   [15:0] Y0_4xDP;
  wire   [15:0] Y1_0xDP;
  wire   [15:0] Y1_1xDP;
  wire   [15:0] Y1_2xDP;
  wire   [15:0] Y1_3xDP;
  wire   [15:0] Y1_4xDP;
  wire   [15:0] Y0xorY12xD;
  wire   [11:0] Y0xorY1xD;
  wire   [15:0] Y0mulY1xD;
  wire   [31:0] InvUnmappedxD;
  wire   [15:0] InverterOutxD;
  wire   [63:0] mul_y0y1_FFxDN;
  wire   [7:0] inverter_gf24_AmulBxD;
  wire   [7:0] inverter_gf24_ExD;
  wire   [7:0] inverter_gf24_pipelinedBxDP;
  wire   [7:0] inverter_gf24_pipelinedAxDP;
  wire   [7:0] inverter_gf24_BxDP;
  wire   [7:0] inverter_gf24_AxDP;
  wire   [31:0] inverter_gf24_a_mul_b_FFxDN;
  wire   [31:0] inverter_gf24_a_mul_e_FFxDN;
  wire   [31:0] inverter_gf24_b_mul_e_FFxDN;
  wire   [63:0] mult_msb_FFxDN;
  wire   [63:0] mult_lsb_FFxDN;

  DFF_X1 mappedxDP_reg_3__7_ ( .D(mappedxD_3__7_), .CK(ClkxCI), .Q(Y1xD[15]), 
        .QN(n42) );
  DFF_X1 mappedxDP_reg_3__6_ ( .D(mappedxD_3__6_), .CK(ClkxCI), .Q(Y1xD[14]), 
        .QN(n44) );
  DFF_X1 mappedxDP_reg_3__5_ ( .D(mappedxD_3__5_), .CK(ClkxCI), .Q(Y1xD[13]), 
        .QN(n46) );
  DFF_X1 mappedxDP_reg_3__4_ ( .D(mappedxD_3__4_), .CK(ClkxCI), .Q(Y1xD[12]), 
        .QN(n48) );
  DFF_X1 mappedxDP_reg_3__3_ ( .D(mappedxD_3__3_), .CK(ClkxCI), .Q(Y0xD[15]), 
        .QN(n41) );
  DFF_X1 mappedxDP_reg_3__2_ ( .D(XxDI[24]), .CK(ClkxCI), .Q(Y0xD[14]), .QN(
        n43) );
  DFF_X1 mappedxDP_reg_3__1_ ( .D(mappedxD_3__1_), .CK(ClkxCI), .Q(Y0xD[13]), 
        .QN(n45) );
  DFF_X1 mappedxDP_reg_3__0_ ( .D(mappedxD_3__0_), .CK(ClkxCI), .Q(Y0xD[12]), 
        .QN(n47) );
  DFF_X1 mappedxDP_reg_2__7_ ( .D(mappedxD_2__7_), .CK(ClkxCI), .Q(Y1xD[11]), 
        .QN(n50) );
  DFF_X1 mappedxDP_reg_2__6_ ( .D(mappedxD_2__6_), .CK(ClkxCI), .Q(Y1xD[10]), 
        .QN(n52) );
  DFF_X1 mappedxDP_reg_2__5_ ( .D(mappedxD_2__5_), .CK(ClkxCI), .Q(Y1xD[9]), 
        .QN(n54) );
  DFF_X1 mappedxDP_reg_2__4_ ( .D(mappedxD_2__4_), .CK(ClkxCI), .Q(Y1xD[8]), 
        .QN(n56) );
  DFF_X1 mappedxDP_reg_2__3_ ( .D(mappedxD_2__3_), .CK(ClkxCI), .Q(Y0xD[11]), 
        .QN(n49) );
  DFF_X1 mappedxDP_reg_2__2_ ( .D(XxDI[16]), .CK(ClkxCI), .Q(Y0xD[10]), .QN(
        n51) );
  DFF_X1 mappedxDP_reg_2__1_ ( .D(mappedxD_2__1_), .CK(ClkxCI), .Q(Y0xD[9]), 
        .QN(n53) );
  DFF_X1 mappedxDP_reg_2__0_ ( .D(mappedxD_2__0_), .CK(ClkxCI), .Q(Y0xD[8]), 
        .QN(n55) );
  DFF_X1 mappedxDP_reg_1__7_ ( .D(mappedxD_1__7_), .CK(ClkxCI), .Q(Y1xD[7]), 
        .QN(n58) );
  DFF_X1 mappedxDP_reg_1__6_ ( .D(mappedxD_1__6_), .CK(ClkxCI), .Q(Y1xD[6]), 
        .QN(n60) );
  DFF_X1 mappedxDP_reg_1__5_ ( .D(mappedxD_1__5_), .CK(ClkxCI), .Q(Y1xD[5]), 
        .QN(n62) );
  DFF_X1 mappedxDP_reg_1__4_ ( .D(mappedxD_1__4_), .CK(ClkxCI), .Q(Y1xD[4]), 
        .QN(n64) );
  DFF_X1 mappedxDP_reg_1__3_ ( .D(mappedxD_1__3_), .CK(ClkxCI), .Q(Y0xD[7]), 
        .QN(n57) );
  DFF_X1 mappedxDP_reg_1__2_ ( .D(XxDI[8]), .CK(ClkxCI), .Q(Y0xD[6]), .QN(n59)
         );
  DFF_X1 mappedxDP_reg_1__1_ ( .D(mappedxD_1__1_), .CK(ClkxCI), .Q(Y0xD[5]), 
        .QN(n61) );
  DFF_X1 mappedxDP_reg_1__0_ ( .D(mappedxD_1__0_), .CK(ClkxCI), .Q(Y0xD[4]), 
        .QN(n63) );
  DFF_X1 mappedxDP_reg_0__7_ ( .D(mappedxD_0__7_), .CK(ClkxCI), .Q(Y1xD[3]), 
        .QN(n66) );
  DFF_X1 mappedxDP_reg_0__6_ ( .D(mappedxD_0__6_), .CK(ClkxCI), .Q(Y1xD[2]), 
        .QN(n68) );
  DFF_X1 mappedxDP_reg_0__5_ ( .D(mappedxD_0__5_), .CK(ClkxCI), .Q(Y1xD[1]), 
        .QN(n70) );
  DFF_X1 mappedxDP_reg_0__4_ ( .D(mappedxD_0__4_), .CK(ClkxCI), .Q(Y1xD[0]), 
        .QN(n72) );
  DFF_X1 mappedxDP_reg_0__3_ ( .D(mappedxD_0__3_), .CK(ClkxCI), .Q(Y0xD[3]), 
        .QN(n65) );
  DFF_X1 mappedxDP_reg_0__2_ ( .D(XxDI[0]), .CK(ClkxCI), .Q(Y0xD[2]), .QN(n67)
         );
  DFF_X1 mappedxDP_reg_0__1_ ( .D(mappedxD_0__1_), .CK(ClkxCI), .Q(Y0xD[1]), 
        .QN(n69) );
  DFF_X1 mappedxDP_reg_0__0_ ( .D(mappedxD_0__0_), .CK(ClkxCI), .Q(Y0xD[0]), 
        .QN(n71) );
  DFF_X1 Y0xorY12xDP_reg_3__3_ ( .D(Y0xorY12xD[15]), .CK(ClkxCI), .Q(), .QN(
        n73) );
  DFF_X1 InverterInxDP_reg_3__3_ ( .D(InverterInxD[15]), .CK(ClkxCI), .Q(
        InverterInxDP[15]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_3__2_ ( .D(Y0xorY12xD[14]), .CK(ClkxCI), .Q(), .QN(
        n74) );
  DFF_X1 InverterInxDP_reg_3__2_ ( .D(InverterInxD[14]), .CK(ClkxCI), .Q(
        InverterInxDP[14]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_3__1_ ( .D(Y0xorY12xD[13]), .CK(ClkxCI), .Q(), .QN(
        n75) );
  DFF_X1 InverterInxDP_reg_3__1_ ( .D(InverterInxD[13]), .CK(ClkxCI), .Q(
        InverterInxDP[13]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_3__0_ ( .D(Y0xorY12xD[12]), .CK(ClkxCI), .Q(), .QN(
        n76) );
  DFF_X1 InverterInxDP_reg_3__0_ ( .D(InverterInxD[12]), .CK(ClkxCI), .Q(
        InverterInxDP[12]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_2__3_ ( .D(Y0xorY12xD[11]), .CK(ClkxCI), .Q(), .QN(
        n77) );
  DFF_X1 InverterInxDP_reg_2__3_ ( .D(InverterInxD[11]), .CK(ClkxCI), .Q(
        InverterInxDP[11]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_2__2_ ( .D(Y0xorY12xD[10]), .CK(ClkxCI), .Q(), .QN(
        n78) );
  DFF_X1 InverterInxDP_reg_2__2_ ( .D(InverterInxD[10]), .CK(ClkxCI), .Q(
        InverterInxDP[10]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_2__1_ ( .D(Y0xorY12xD[9]), .CK(ClkxCI), .Q(), .QN(n79) );
  DFF_X1 InverterInxDP_reg_2__1_ ( .D(InverterInxD[9]), .CK(ClkxCI), .Q(
        InverterInxDP[9]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_2__0_ ( .D(Y0xorY12xD[8]), .CK(ClkxCI), .Q(), .QN(n80) );
  DFF_X1 InverterInxDP_reg_2__0_ ( .D(InverterInxD[8]), .CK(ClkxCI), .Q(
        InverterInxDP[8]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_1__3_ ( .D(Y0xorY12xD[7]), .CK(ClkxCI), .Q(), .QN(n81) );
  DFF_X1 InverterInxDP_reg_1__3_ ( .D(InverterInxD[7]), .CK(ClkxCI), .Q(
        InverterInxDP[7]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_1__2_ ( .D(Y0xorY12xD[6]), .CK(ClkxCI), .Q(), .QN(n82) );
  DFF_X1 InverterInxDP_reg_1__2_ ( .D(InverterInxD[6]), .CK(ClkxCI), .Q(
        InverterInxDP[6]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_1__1_ ( .D(Y0xorY12xD[5]), .CK(ClkxCI), .Q(), .QN(n83) );
  DFF_X1 InverterInxDP_reg_1__1_ ( .D(InverterInxD[5]), .CK(ClkxCI), .Q(
        InverterInxDP[5]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_1__0_ ( .D(Y0xorY12xD[4]), .CK(ClkxCI), .Q(), .QN(n84) );
  DFF_X1 InverterInxDP_reg_1__0_ ( .D(InverterInxD[4]), .CK(ClkxCI), .Q(
        InverterInxDP[4]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_0__3_ ( .D(Y0xorY12xD[3]), .CK(ClkxCI), .Q(), .QN(n85) );
  DFF_X1 InverterInxDP_reg_0__3_ ( .D(InverterInxD[3]), .CK(ClkxCI), .Q(
        InverterInxDP[3]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_0__2_ ( .D(Y0xorY12xD[2]), .CK(ClkxCI), .Q(), .QN(n86) );
  DFF_X1 InverterInxDP_reg_0__2_ ( .D(InverterInxD[2]), .CK(ClkxCI), .Q(
        InverterInxDP[2]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_0__1_ ( .D(Y0xorY12xD[1]), .CK(ClkxCI), .Q(), .QN(n87) );
  DFF_X1 InverterInxDP_reg_0__1_ ( .D(InverterInxD[1]), .CK(ClkxCI), .Q(
        InverterInxDP[1]), .QN() );
  DFF_X1 Y0xorY12xDP_reg_0__0_ ( .D(Y0xorY12xD[0]), .CK(ClkxCI), .Q(), .QN(n88) );
  DFF_X1 InverterInxDP_reg_0__0_ ( .D(InverterInxD[0]), .CK(ClkxCI), .Q(
        InverterInxDP[0]), .QN() );
  DFF_X1 Y0_0xDP_reg_3__3_ ( .D(Y0xD[15]), .CK(ClkxCI), .Q(Y0_0xDP[15]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_3__2_ ( .D(Y0xD[14]), .CK(ClkxCI), .Q(Y0_0xDP[14]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_3__1_ ( .D(Y0xD[13]), .CK(ClkxCI), .Q(Y0_0xDP[13]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_3__0_ ( .D(Y0xD[12]), .CK(ClkxCI), .Q(Y0_0xDP[12]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_2__3_ ( .D(Y0xD[11]), .CK(ClkxCI), .Q(Y0_0xDP[11]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_2__2_ ( .D(Y0xD[10]), .CK(ClkxCI), .Q(Y0_0xDP[10]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_2__1_ ( .D(Y0xD[9]), .CK(ClkxCI), .Q(Y0_0xDP[9]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_2__0_ ( .D(Y0xD[8]), .CK(ClkxCI), .Q(Y0_0xDP[8]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_1__3_ ( .D(Y0xD[7]), .CK(ClkxCI), .Q(Y0_0xDP[7]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_1__2_ ( .D(Y0xD[6]), .CK(ClkxCI), .Q(Y0_0xDP[6]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_1__1_ ( .D(Y0xD[5]), .CK(ClkxCI), .Q(Y0_0xDP[5]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_1__0_ ( .D(Y0xD[4]), .CK(ClkxCI), .Q(Y0_0xDP[4]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_0__3_ ( .D(Y0xD[3]), .CK(ClkxCI), .Q(Y0_0xDP[3]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_0__2_ ( .D(Y0xD[2]), .CK(ClkxCI), .Q(Y0_0xDP[2]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_0__1_ ( .D(Y0xD[1]), .CK(ClkxCI), .Q(Y0_0xDP[1]), .QN()
         );
  DFF_X1 Y0_0xDP_reg_0__0_ ( .D(Y0xD[0]), .CK(ClkxCI), .Q(Y0_0xDP[0]), .QN()
         );
  DFF_X1 Y0_1xDP_reg_3__3_ ( .D(Y0_0xDP[15]), .CK(ClkxCI), .Q(Y0_1xDP[15]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_3__2_ ( .D(Y0_0xDP[14]), .CK(ClkxCI), .Q(Y0_1xDP[14]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_3__1_ ( .D(Y0_0xDP[13]), .CK(ClkxCI), .Q(Y0_1xDP[13]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_3__0_ ( .D(Y0_0xDP[12]), .CK(ClkxCI), .Q(Y0_1xDP[12]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_2__3_ ( .D(Y0_0xDP[11]), .CK(ClkxCI), .Q(Y0_1xDP[11]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_2__2_ ( .D(Y0_0xDP[10]), .CK(ClkxCI), .Q(Y0_1xDP[10]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_2__1_ ( .D(Y0_0xDP[9]), .CK(ClkxCI), .Q(Y0_1xDP[9]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_2__0_ ( .D(Y0_0xDP[8]), .CK(ClkxCI), .Q(Y0_1xDP[8]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_1__3_ ( .D(Y0_0xDP[7]), .CK(ClkxCI), .Q(Y0_1xDP[7]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_1__2_ ( .D(Y0_0xDP[6]), .CK(ClkxCI), .Q(Y0_1xDP[6]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_1__1_ ( .D(Y0_0xDP[5]), .CK(ClkxCI), .Q(Y0_1xDP[5]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_1__0_ ( .D(Y0_0xDP[4]), .CK(ClkxCI), .Q(Y0_1xDP[4]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_0__3_ ( .D(Y0_0xDP[3]), .CK(ClkxCI), .Q(Y0_1xDP[3]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_0__2_ ( .D(Y0_0xDP[2]), .CK(ClkxCI), .Q(Y0_1xDP[2]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_0__1_ ( .D(Y0_0xDP[1]), .CK(ClkxCI), .Q(Y0_1xDP[1]), 
        .QN() );
  DFF_X1 Y0_1xDP_reg_0__0_ ( .D(Y0_0xDP[0]), .CK(ClkxCI), .Q(Y0_1xDP[0]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_3__3_ ( .D(Y0_1xDP[15]), .CK(ClkxCI), .Q(Y0_2xDP[15]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_3__2_ ( .D(Y0_1xDP[14]), .CK(ClkxCI), .Q(Y0_2xDP[14]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_3__1_ ( .D(Y0_1xDP[13]), .CK(ClkxCI), .Q(Y0_2xDP[13]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_3__0_ ( .D(Y0_1xDP[12]), .CK(ClkxCI), .Q(Y0_2xDP[12]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_2__3_ ( .D(Y0_1xDP[11]), .CK(ClkxCI), .Q(Y0_2xDP[11]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_2__2_ ( .D(Y0_1xDP[10]), .CK(ClkxCI), .Q(Y0_2xDP[10]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_2__1_ ( .D(Y0_1xDP[9]), .CK(ClkxCI), .Q(Y0_2xDP[9]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_2__0_ ( .D(Y0_1xDP[8]), .CK(ClkxCI), .Q(Y0_2xDP[8]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_1__3_ ( .D(Y0_1xDP[7]), .CK(ClkxCI), .Q(Y0_2xDP[7]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_1__2_ ( .D(Y0_1xDP[6]), .CK(ClkxCI), .Q(Y0_2xDP[6]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_1__1_ ( .D(Y0_1xDP[5]), .CK(ClkxCI), .Q(Y0_2xDP[5]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_1__0_ ( .D(Y0_1xDP[4]), .CK(ClkxCI), .Q(Y0_2xDP[4]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_0__3_ ( .D(Y0_1xDP[3]), .CK(ClkxCI), .Q(Y0_2xDP[3]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_0__2_ ( .D(Y0_1xDP[2]), .CK(ClkxCI), .Q(Y0_2xDP[2]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_0__1_ ( .D(Y0_1xDP[1]), .CK(ClkxCI), .Q(Y0_2xDP[1]), 
        .QN() );
  DFF_X1 Y0_2xDP_reg_0__0_ ( .D(Y0_1xDP[0]), .CK(ClkxCI), .Q(Y0_2xDP[0]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_3__3_ ( .D(Y0_2xDP[15]), .CK(ClkxCI), .Q(Y0_3xDP[15]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_3__2_ ( .D(Y0_2xDP[14]), .CK(ClkxCI), .Q(Y0_3xDP[14]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_3__1_ ( .D(Y0_2xDP[13]), .CK(ClkxCI), .Q(Y0_3xDP[13]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_3__0_ ( .D(Y0_2xDP[12]), .CK(ClkxCI), .Q(Y0_3xDP[12]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_2__3_ ( .D(Y0_2xDP[11]), .CK(ClkxCI), .Q(Y0_3xDP[11]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_2__2_ ( .D(Y0_2xDP[10]), .CK(ClkxCI), .Q(Y0_3xDP[10]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_2__1_ ( .D(Y0_2xDP[9]), .CK(ClkxCI), .Q(Y0_3xDP[9]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_2__0_ ( .D(Y0_2xDP[8]), .CK(ClkxCI), .Q(Y0_3xDP[8]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_1__3_ ( .D(Y0_2xDP[7]), .CK(ClkxCI), .Q(Y0_3xDP[7]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_1__2_ ( .D(Y0_2xDP[6]), .CK(ClkxCI), .Q(Y0_3xDP[6]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_1__1_ ( .D(Y0_2xDP[5]), .CK(ClkxCI), .Q(Y0_3xDP[5]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_1__0_ ( .D(Y0_2xDP[4]), .CK(ClkxCI), .Q(Y0_3xDP[4]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_0__3_ ( .D(Y0_2xDP[3]), .CK(ClkxCI), .Q(Y0_3xDP[3]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_0__2_ ( .D(Y0_2xDP[2]), .CK(ClkxCI), .Q(Y0_3xDP[2]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_0__1_ ( .D(Y0_2xDP[1]), .CK(ClkxCI), .Q(Y0_3xDP[1]), 
        .QN() );
  DFF_X1 Y0_3xDP_reg_0__0_ ( .D(Y0_2xDP[0]), .CK(ClkxCI), .Q(Y0_3xDP[0]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_3__3_ ( .D(Y0_3xDP[15]), .CK(ClkxCI), .Q(Y0_4xDP[15]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_3__2_ ( .D(Y0_3xDP[14]), .CK(ClkxCI), .Q(Y0_4xDP[14]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_3__1_ ( .D(Y0_3xDP[13]), .CK(ClkxCI), .Q(Y0_4xDP[13]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_3__0_ ( .D(Y0_3xDP[12]), .CK(ClkxCI), .Q(Y0_4xDP[12]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_2__3_ ( .D(Y0_3xDP[11]), .CK(ClkxCI), .Q(Y0_4xDP[11]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_2__2_ ( .D(Y0_3xDP[10]), .CK(ClkxCI), .Q(Y0_4xDP[10]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_2__1_ ( .D(Y0_3xDP[9]), .CK(ClkxCI), .Q(Y0_4xDP[9]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_2__0_ ( .D(Y0_3xDP[8]), .CK(ClkxCI), .Q(Y0_4xDP[8]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_1__3_ ( .D(Y0_3xDP[7]), .CK(ClkxCI), .Q(Y0_4xDP[7]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_1__2_ ( .D(Y0_3xDP[6]), .CK(ClkxCI), .Q(Y0_4xDP[6]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_1__1_ ( .D(Y0_3xDP[5]), .CK(ClkxCI), .Q(Y0_4xDP[5]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_1__0_ ( .D(Y0_3xDP[4]), .CK(ClkxCI), .Q(Y0_4xDP[4]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_0__3_ ( .D(Y0_3xDP[3]), .CK(ClkxCI), .Q(Y0_4xDP[3]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_0__2_ ( .D(Y0_3xDP[2]), .CK(ClkxCI), .Q(Y0_4xDP[2]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_0__1_ ( .D(Y0_3xDP[1]), .CK(ClkxCI), .Q(Y0_4xDP[1]), 
        .QN() );
  DFF_X1 Y0_4xDP_reg_0__0_ ( .D(Y0_3xDP[0]), .CK(ClkxCI), .Q(Y0_4xDP[0]), 
        .QN() );
  DFF_X1 Y1_0xDP_reg_3__3_ ( .D(Y1xD[15]), .CK(ClkxCI), .Q(Y1_0xDP[15]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_3__2_ ( .D(Y1xD[14]), .CK(ClkxCI), .Q(Y1_0xDP[14]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_3__1_ ( .D(Y1xD[13]), .CK(ClkxCI), .Q(Y1_0xDP[13]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_3__0_ ( .D(Y1xD[12]), .CK(ClkxCI), .Q(Y1_0xDP[12]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_2__3_ ( .D(Y1xD[11]), .CK(ClkxCI), .Q(Y1_0xDP[11]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_2__2_ ( .D(Y1xD[10]), .CK(ClkxCI), .Q(Y1_0xDP[10]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_2__1_ ( .D(Y1xD[9]), .CK(ClkxCI), .Q(Y1_0xDP[9]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_2__0_ ( .D(Y1xD[8]), .CK(ClkxCI), .Q(Y1_0xDP[8]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_1__3_ ( .D(Y1xD[7]), .CK(ClkxCI), .Q(Y1_0xDP[7]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_1__2_ ( .D(Y1xD[6]), .CK(ClkxCI), .Q(Y1_0xDP[6]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_1__1_ ( .D(Y1xD[5]), .CK(ClkxCI), .Q(Y1_0xDP[5]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_1__0_ ( .D(Y1xD[4]), .CK(ClkxCI), .Q(Y1_0xDP[4]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_0__3_ ( .D(Y1xD[3]), .CK(ClkxCI), .Q(Y1_0xDP[3]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_0__2_ ( .D(Y1xD[2]), .CK(ClkxCI), .Q(Y1_0xDP[2]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_0__1_ ( .D(Y1xD[1]), .CK(ClkxCI), .Q(Y1_0xDP[1]), .QN()
         );
  DFF_X1 Y1_0xDP_reg_0__0_ ( .D(Y1xD[0]), .CK(ClkxCI), .Q(Y1_0xDP[0]), .QN()
         );
  DFF_X1 Y1_1xDP_reg_3__3_ ( .D(Y1_0xDP[15]), .CK(ClkxCI), .Q(Y1_1xDP[15]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_3__2_ ( .D(Y1_0xDP[14]), .CK(ClkxCI), .Q(Y1_1xDP[14]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_3__1_ ( .D(Y1_0xDP[13]), .CK(ClkxCI), .Q(Y1_1xDP[13]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_3__0_ ( .D(Y1_0xDP[12]), .CK(ClkxCI), .Q(Y1_1xDP[12]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_2__3_ ( .D(Y1_0xDP[11]), .CK(ClkxCI), .Q(Y1_1xDP[11]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_2__2_ ( .D(Y1_0xDP[10]), .CK(ClkxCI), .Q(Y1_1xDP[10]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_2__1_ ( .D(Y1_0xDP[9]), .CK(ClkxCI), .Q(Y1_1xDP[9]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_2__0_ ( .D(Y1_0xDP[8]), .CK(ClkxCI), .Q(Y1_1xDP[8]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_1__3_ ( .D(Y1_0xDP[7]), .CK(ClkxCI), .Q(Y1_1xDP[7]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_1__2_ ( .D(Y1_0xDP[6]), .CK(ClkxCI), .Q(Y1_1xDP[6]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_1__1_ ( .D(Y1_0xDP[5]), .CK(ClkxCI), .Q(Y1_1xDP[5]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_1__0_ ( .D(Y1_0xDP[4]), .CK(ClkxCI), .Q(Y1_1xDP[4]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_0__3_ ( .D(Y1_0xDP[3]), .CK(ClkxCI), .Q(Y1_1xDP[3]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_0__2_ ( .D(Y1_0xDP[2]), .CK(ClkxCI), .Q(Y1_1xDP[2]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_0__1_ ( .D(Y1_0xDP[1]), .CK(ClkxCI), .Q(Y1_1xDP[1]), 
        .QN() );
  DFF_X1 Y1_1xDP_reg_0__0_ ( .D(Y1_0xDP[0]), .CK(ClkxCI), .Q(Y1_1xDP[0]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_3__3_ ( .D(Y1_1xDP[15]), .CK(ClkxCI), .Q(Y1_2xDP[15]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_3__2_ ( .D(Y1_1xDP[14]), .CK(ClkxCI), .Q(Y1_2xDP[14]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_3__1_ ( .D(Y1_1xDP[13]), .CK(ClkxCI), .Q(Y1_2xDP[13]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_3__0_ ( .D(Y1_1xDP[12]), .CK(ClkxCI), .Q(Y1_2xDP[12]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_2__3_ ( .D(Y1_1xDP[11]), .CK(ClkxCI), .Q(Y1_2xDP[11]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_2__2_ ( .D(Y1_1xDP[10]), .CK(ClkxCI), .Q(Y1_2xDP[10]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_2__1_ ( .D(Y1_1xDP[9]), .CK(ClkxCI), .Q(Y1_2xDP[9]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_2__0_ ( .D(Y1_1xDP[8]), .CK(ClkxCI), .Q(Y1_2xDP[8]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_1__3_ ( .D(Y1_1xDP[7]), .CK(ClkxCI), .Q(Y1_2xDP[7]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_1__2_ ( .D(Y1_1xDP[6]), .CK(ClkxCI), .Q(Y1_2xDP[6]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_1__1_ ( .D(Y1_1xDP[5]), .CK(ClkxCI), .Q(Y1_2xDP[5]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_1__0_ ( .D(Y1_1xDP[4]), .CK(ClkxCI), .Q(Y1_2xDP[4]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_0__3_ ( .D(Y1_1xDP[3]), .CK(ClkxCI), .Q(Y1_2xDP[3]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_0__2_ ( .D(Y1_1xDP[2]), .CK(ClkxCI), .Q(Y1_2xDP[2]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_0__1_ ( .D(Y1_1xDP[1]), .CK(ClkxCI), .Q(Y1_2xDP[1]), 
        .QN() );
  DFF_X1 Y1_2xDP_reg_0__0_ ( .D(Y1_1xDP[0]), .CK(ClkxCI), .Q(Y1_2xDP[0]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_3__3_ ( .D(Y1_2xDP[15]), .CK(ClkxCI), .Q(Y1_3xDP[15]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_3__3_ ( .D(Y1_3xDP[15]), .CK(ClkxCI), .Q(Y1_4xDP[15]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_3__2_ ( .D(Y1_2xDP[14]), .CK(ClkxCI), .Q(Y1_3xDP[14]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_3__2_ ( .D(Y1_3xDP[14]), .CK(ClkxCI), .Q(Y1_4xDP[14]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_3__1_ ( .D(Y1_2xDP[13]), .CK(ClkxCI), .Q(Y1_3xDP[13]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_3__1_ ( .D(Y1_3xDP[13]), .CK(ClkxCI), .Q(Y1_4xDP[13]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_3__0_ ( .D(Y1_2xDP[12]), .CK(ClkxCI), .Q(Y1_3xDP[12]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_3__0_ ( .D(Y1_3xDP[12]), .CK(ClkxCI), .Q(Y1_4xDP[12]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_2__3_ ( .D(Y1_2xDP[11]), .CK(ClkxCI), .Q(Y1_3xDP[11]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_2__3_ ( .D(Y1_3xDP[11]), .CK(ClkxCI), .Q(Y1_4xDP[11]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_2__2_ ( .D(Y1_2xDP[10]), .CK(ClkxCI), .Q(Y1_3xDP[10]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_2__2_ ( .D(Y1_3xDP[10]), .CK(ClkxCI), .Q(Y1_4xDP[10]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_2__1_ ( .D(Y1_2xDP[9]), .CK(ClkxCI), .Q(Y1_3xDP[9]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_2__1_ ( .D(Y1_3xDP[9]), .CK(ClkxCI), .Q(Y1_4xDP[9]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_2__0_ ( .D(Y1_2xDP[8]), .CK(ClkxCI), .Q(Y1_3xDP[8]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_2__0_ ( .D(Y1_3xDP[8]), .CK(ClkxCI), .Q(Y1_4xDP[8]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_1__3_ ( .D(Y1_2xDP[7]), .CK(ClkxCI), .Q(Y1_3xDP[7]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_1__3_ ( .D(Y1_3xDP[7]), .CK(ClkxCI), .Q(Y1_4xDP[7]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_1__2_ ( .D(Y1_2xDP[6]), .CK(ClkxCI), .Q(Y1_3xDP[6]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_1__2_ ( .D(Y1_3xDP[6]), .CK(ClkxCI), .Q(Y1_4xDP[6]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_1__1_ ( .D(Y1_2xDP[5]), .CK(ClkxCI), .Q(Y1_3xDP[5]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_1__1_ ( .D(Y1_3xDP[5]), .CK(ClkxCI), .Q(Y1_4xDP[5]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_1__0_ ( .D(Y1_2xDP[4]), .CK(ClkxCI), .Q(Y1_3xDP[4]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_1__0_ ( .D(Y1_3xDP[4]), .CK(ClkxCI), .Q(Y1_4xDP[4]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_0__3_ ( .D(Y1_2xDP[3]), .CK(ClkxCI), .Q(Y1_3xDP[3]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_0__3_ ( .D(Y1_3xDP[3]), .CK(ClkxCI), .Q(Y1_4xDP[3]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_0__2_ ( .D(Y1_2xDP[2]), .CK(ClkxCI), .Q(Y1_3xDP[2]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_0__2_ ( .D(Y1_3xDP[2]), .CK(ClkxCI), .Q(Y1_4xDP[2]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_0__1_ ( .D(Y1_2xDP[1]), .CK(ClkxCI), .Q(Y1_3xDP[1]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_0__1_ ( .D(Y1_3xDP[1]), .CK(ClkxCI), .Q(Y1_4xDP[1]), 
        .QN() );
  DFF_X1 Y1_3xDP_reg_0__0_ ( .D(Y1_2xDP[0]), .CK(ClkxCI), .Q(Y1_3xDP[0]), 
        .QN() );
  DFF_X1 Y1_4xDP_reg_0__0_ ( .D(Y1_3xDP[0]), .CK(ClkxCI), .Q(Y1_4xDP[0]), 
        .QN() );
  INV_X2 U75 ( .A(n92), .ZN(n91) );
  INV_X2 U76 ( .A(n100), .ZN(n99) );
  INV_X2 U77 ( .A(n108), .ZN(n107) );
  INV_X2 U78 ( .A(n116), .ZN(n115) );
  INV_X2 U79 ( .A(n94), .ZN(n93) );
  INV_X2 U80 ( .A(n102), .ZN(n101) );
  INV_X2 U81 ( .A(n110), .ZN(n109) );
  INV_X2 U82 ( .A(n118), .ZN(n117) );
  INV_X2 U83 ( .A(n114), .ZN(n113) );
  INV_X2 U84 ( .A(n106), .ZN(n105) );
  INV_X2 U85 ( .A(n98), .ZN(n97) );
  INV_X2 U86 ( .A(n90), .ZN(n89) );
  INV_X2 U87 ( .A(n120), .ZN(n119) );
  INV_X2 U88 ( .A(n112), .ZN(n111) );
  INV_X2 U89 ( .A(n104), .ZN(n103) );
  INV_X2 U90 ( .A(n96), .ZN(n95) );
  INV_X1 U91 ( .A(InverterOutxD[0]), .ZN(n90) );
  INV_X1 U92 ( .A(InverterOutxD[1]), .ZN(n92) );
  INV_X1 U93 ( .A(InverterOutxD[2]), .ZN(n94) );
  INV_X1 U94 ( .A(InverterOutxD[3]), .ZN(n96) );
  INV_X1 U95 ( .A(InverterOutxD[4]), .ZN(n98) );
  INV_X1 U96 ( .A(InverterOutxD[5]), .ZN(n100) );
  INV_X1 U97 ( .A(InverterOutxD[6]), .ZN(n102) );
  INV_X1 U98 ( .A(InverterOutxD[7]), .ZN(n104) );
  INV_X1 U99 ( .A(InverterOutxD[8]), .ZN(n106) );
  INV_X1 U100 ( .A(InverterOutxD[9]), .ZN(n108) );
  INV_X1 U101 ( .A(InverterOutxD[10]), .ZN(n110) );
  INV_X1 U102 ( .A(InverterOutxD[11]), .ZN(n112) );
  INV_X1 U103 ( .A(InverterOutxD[12]), .ZN(n114) );
  INV_X1 U104 ( .A(InverterOutxD[13]), .ZN(n116) );
  INV_X1 U105 ( .A(InverterOutxD[14]), .ZN(n118) );
  INV_X1 U106 ( .A(InverterOutxD[15]), .ZN(n120) );
  XNOR2_X1 U108 ( .A(Y0mulY1xD[0]), .B(n88), .ZN(InverterInxD[0]) );
  XNOR2_X1 U109 ( .A(Y0mulY1xD[1]), .B(n87), .ZN(InverterInxD[1]) );
  XNOR2_X1 U110 ( .A(Y0mulY1xD[2]), .B(n86), .ZN(InverterInxD[2]) );
  XNOR2_X1 U111 ( .A(Y0mulY1xD[3]), .B(n85), .ZN(InverterInxD[3]) );
  XNOR2_X1 U112 ( .A(Y0mulY1xD[4]), .B(n84), .ZN(InverterInxD[4]) );
  XNOR2_X1 U113 ( .A(Y0mulY1xD[5]), .B(n83), .ZN(InverterInxD[5]) );
  XNOR2_X1 U114 ( .A(Y0mulY1xD[6]), .B(n82), .ZN(InverterInxD[6]) );
  XNOR2_X1 U115 ( .A(Y0mulY1xD[7]), .B(n81), .ZN(InverterInxD[7]) );
  XNOR2_X1 U116 ( .A(Y0mulY1xD[8]), .B(n80), .ZN(InverterInxD[8]) );
  XNOR2_X1 U117 ( .A(Y0mulY1xD[9]), .B(n79), .ZN(InverterInxD[9]) );
  XNOR2_X1 U118 ( .A(Y0mulY1xD[10]), .B(n78), .ZN(InverterInxD[10]) );
  XNOR2_X1 U119 ( .A(Y0mulY1xD[11]), .B(n77), .ZN(InverterInxD[11]) );
  XNOR2_X1 U120 ( .A(Y0mulY1xD[12]), .B(n76), .ZN(InverterInxD[12]) );
  XNOR2_X1 U121 ( .A(Y0mulY1xD[13]), .B(n75), .ZN(InverterInxD[13]) );
  XNOR2_X1 U122 ( .A(Y0mulY1xD[14]), .B(n74), .ZN(InverterInxD[14]) );
  XNOR2_X1 U123 ( .A(Y0mulY1xD[15]), .B(n73), .ZN(InverterInxD[15]) );
  XOR2_X1 U124 ( .A(n72), .B(n71), .Z(Y0xorY12xD[0]) );
  XOR2_X1 U125 ( .A(n70), .B(n69), .Z(Y0xorY1xD[0]) );
  XOR2_X1 U126 ( .A(n68), .B(n67), .Z(Y0xorY1xD[1]) );
  XOR2_X1 U127 ( .A(n66), .B(n65), .Z(Y0xorY1xD[2]) );
  XOR2_X1 U128 ( .A(n64), .B(n63), .Z(Y0xorY12xD[4]) );
  XOR2_X1 U129 ( .A(n62), .B(n61), .Z(Y0xorY1xD[3]) );
  XOR2_X1 U130 ( .A(n60), .B(n59), .Z(Y0xorY1xD[4]) );
  XOR2_X1 U131 ( .A(n58), .B(n57), .Z(Y0xorY1xD[5]) );
  XOR2_X1 U132 ( .A(n56), .B(n55), .Z(Y0xorY12xD[8]) );
  XOR2_X1 U133 ( .A(n54), .B(n53), .Z(Y0xorY1xD[6]) );
  XOR2_X1 U134 ( .A(n52), .B(n51), .Z(Y0xorY1xD[7]) );
  XOR2_X1 U135 ( .A(n50), .B(n49), .Z(Y0xorY1xD[8]) );
  XOR2_X1 U136 ( .A(n48), .B(n47), .Z(Y0xorY12xD[12]) );
  XOR2_X1 U137 ( .A(n46), .B(n45), .Z(Y0xorY1xD[9]) );
  XOR2_X1 U138 ( .A(n44), .B(n43), .Z(Y0xorY1xD[10]) );
  XOR2_X1 U139 ( .A(n42), .B(n41), .Z(Y0xorY1xD[11]) );
  INV_X1 U140 ( .A(InvMappedxD_0__6_), .ZN(QxDO[6]) );
  INV_X1 U141 ( .A(InvMappedxD_0__5_), .ZN(QxDO[5]) );
  INV_X1 U142 ( .A(InvMappedxD_0__1_), .ZN(QxDO[1]) );
  INV_X1 U143 ( .A(InvMappedxD_0__0_), .ZN(QxDO[0]) );
  XNOR2_X1 input_mapping_3_U14 ( .A(input_mapping_3_n23), .B(
        input_mapping_3_n22), .ZN(mappedxD_3__7_) );
  XOR2_X1 input_mapping_3_U13 ( .A(XxDI[28]), .B(mappedxD_3__1_), .Z(
        mappedxD_3__6_) );
  XNOR2_X1 input_mapping_3_U12 ( .A(input_mapping_3_n21), .B(
        input_mapping_3_n20), .ZN(mappedxD_3__5_) );
  XNOR2_X1 input_mapping_3_U11 ( .A(XxDI[24]), .B(input_mapping_3_n22), .ZN(
        mappedxD_3__4_) );
  XNOR2_X1 input_mapping_3_U10 ( .A(XxDI[31]), .B(input_mapping_3_n21), .ZN(
        input_mapping_3_n22) );
  XNOR2_X1 input_mapping_3_U9 ( .A(input_mapping_3_n19), .B(
        input_mapping_3_n18), .ZN(mappedxD_3__3_) );
  XNOR2_X1 input_mapping_3_U8 ( .A(input_mapping_3_n20), .B(XxDI[27]), .ZN(
        input_mapping_3_n18) );
  XNOR2_X1 input_mapping_3_U7 ( .A(XxDI[31]), .B(XxDI[28]), .ZN(
        input_mapping_3_n19) );
  XOR2_X1 input_mapping_3_U6 ( .A(XxDI[24]), .B(input_mapping_3_n21), .Z(
        mappedxD_3__1_) );
  XOR2_X1 input_mapping_3_U5 ( .A(XxDI[30]), .B(XxDI[29]), .Z(
        input_mapping_3_n21) );
  XNOR2_X1 input_mapping_3_U4 ( .A(input_mapping_3_n23), .B(
        input_mapping_3_n17), .ZN(mappedxD_3__0_) );
  XNOR2_X1 input_mapping_3_U3 ( .A(XxDI[30]), .B(XxDI[27]), .ZN(
        input_mapping_3_n17) );
  XNOR2_X1 input_mapping_3_U2 ( .A(XxDI[26]), .B(input_mapping_3_n20), .ZN(
        input_mapping_3_n23) );
  XNOR2_X1 input_mapping_3_U1 ( .A(XxDI[24]), .B(XxDI[25]), .ZN(
        input_mapping_3_n20) );
  XOR2_X1 square_scaler_gf24_3_U3 ( .A(Y0xorY12xD[12]), .B(Y0xorY1xD[10]), .Z(
        Y0xorY12xD[15]) );
  XOR2_X1 square_scaler_gf24_3_U2 ( .A(Y0xorY1xD[9]), .B(Y0xorY1xD[11]), .Z(
        Y0xorY12xD[14]) );
  XOR2_X1 square_scaler_gf24_3_U1 ( .A(Y0xorY12xD[12]), .B(Y0xorY1xD[9]), .Z(
        Y0xorY12xD[13]) );
  XOR2_X1 output_mapping_3_U11 ( .A(InvUnmappedxD[27]), .B(InvUnmappedxD[31]), 
        .Z(QxDO[30]) );
  XNOR2_X1 output_mapping_3_U10 ( .A(QxDO[28]), .B(output_mapping_3_n9), .ZN(
        QxDO[27]) );
  XOR2_X1 output_mapping_3_U9 ( .A(QxDO[31]), .B(InvUnmappedxD[31]), .Z(
        QxDO[28]) );
  XNOR2_X1 output_mapping_3_U8 ( .A(output_mapping_3_n8), .B(QxDO[29]), .ZN(
        QxDO[26]) );
  XNOR2_X1 output_mapping_3_U7 ( .A(QxDO[31]), .B(InvUnmappedxD[26]), .ZN(
        output_mapping_3_n8) );
  XOR2_X1 output_mapping_3_U6 ( .A(InvUnmappedxD[30]), .B(InvUnmappedxD[24]), 
        .Z(QxDO[29]) );
  XOR2_X1 output_mapping_3_U5 ( .A(InvUnmappedxD[27]), .B(InvUnmappedxD[29]), 
        .Z(QxDO[31]) );
  XNOR2_X1 output_mapping_3_U4 ( .A(output_mapping_3_n7), .B(InvUnmappedxD[25]), .ZN(QxDO[25]) );
  XNOR2_X1 output_mapping_3_U3 ( .A(InvUnmappedxD[29]), .B(InvUnmappedxD[28]), 
        .ZN(output_mapping_3_n7) );
  XNOR2_X1 output_mapping_3_U2 ( .A(InvUnmappedxD[25]), .B(output_mapping_3_n9), .ZN(QxDO[24]) );
  XNOR2_X1 output_mapping_3_U1 ( .A(InvUnmappedxD[30]), .B(InvUnmappedxD[28]), 
        .ZN(output_mapping_3_n9) );
  XNOR2_X1 input_mapping_2_U14 ( .A(input_mapping_2_n23), .B(
        input_mapping_2_n22), .ZN(mappedxD_2__7_) );
  XOR2_X1 input_mapping_2_U13 ( .A(XxDI[20]), .B(mappedxD_2__1_), .Z(
        mappedxD_2__6_) );
  XNOR2_X1 input_mapping_2_U12 ( .A(input_mapping_2_n21), .B(
        input_mapping_2_n20), .ZN(mappedxD_2__5_) );
  XNOR2_X1 input_mapping_2_U11 ( .A(XxDI[16]), .B(input_mapping_2_n22), .ZN(
        mappedxD_2__4_) );
  XNOR2_X1 input_mapping_2_U10 ( .A(XxDI[23]), .B(input_mapping_2_n21), .ZN(
        input_mapping_2_n22) );
  XNOR2_X1 input_mapping_2_U9 ( .A(input_mapping_2_n19), .B(
        input_mapping_2_n18), .ZN(mappedxD_2__3_) );
  XNOR2_X1 input_mapping_2_U8 ( .A(input_mapping_2_n20), .B(XxDI[19]), .ZN(
        input_mapping_2_n18) );
  XNOR2_X1 input_mapping_2_U7 ( .A(XxDI[23]), .B(XxDI[20]), .ZN(
        input_mapping_2_n19) );
  XOR2_X1 input_mapping_2_U6 ( .A(XxDI[16]), .B(input_mapping_2_n21), .Z(
        mappedxD_2__1_) );
  XOR2_X1 input_mapping_2_U5 ( .A(XxDI[22]), .B(XxDI[21]), .Z(
        input_mapping_2_n21) );
  XNOR2_X1 input_mapping_2_U4 ( .A(input_mapping_2_n23), .B(
        input_mapping_2_n17), .ZN(mappedxD_2__0_) );
  XNOR2_X1 input_mapping_2_U3 ( .A(XxDI[22]), .B(XxDI[19]), .ZN(
        input_mapping_2_n17) );
  XNOR2_X1 input_mapping_2_U2 ( .A(XxDI[18]), .B(input_mapping_2_n20), .ZN(
        input_mapping_2_n23) );
  XNOR2_X1 input_mapping_2_U1 ( .A(XxDI[16]), .B(XxDI[17]), .ZN(
        input_mapping_2_n20) );
  XOR2_X1 square_scaler_gf24_2_U3 ( .A(Y0xorY12xD[8]), .B(Y0xorY1xD[7]), .Z(
        Y0xorY12xD[11]) );
  XOR2_X1 square_scaler_gf24_2_U2 ( .A(Y0xorY1xD[6]), .B(Y0xorY1xD[8]), .Z(
        Y0xorY12xD[10]) );
  XOR2_X1 square_scaler_gf24_2_U1 ( .A(Y0xorY12xD[8]), .B(Y0xorY1xD[6]), .Z(
        Y0xorY12xD[9]) );
  XOR2_X1 output_mapping_2_U11 ( .A(InvUnmappedxD[19]), .B(InvUnmappedxD[23]), 
        .Z(QxDO[22]) );
  XNOR2_X1 output_mapping_2_U10 ( .A(QxDO[20]), .B(output_mapping_2_n9), .ZN(
        QxDO[19]) );
  XOR2_X1 output_mapping_2_U9 ( .A(QxDO[23]), .B(InvUnmappedxD[23]), .Z(
        QxDO[20]) );
  XNOR2_X1 output_mapping_2_U8 ( .A(output_mapping_2_n8), .B(QxDO[21]), .ZN(
        QxDO[18]) );
  XNOR2_X1 output_mapping_2_U7 ( .A(QxDO[23]), .B(InvUnmappedxD[18]), .ZN(
        output_mapping_2_n8) );
  XOR2_X1 output_mapping_2_U6 ( .A(InvUnmappedxD[22]), .B(InvUnmappedxD[16]), 
        .Z(QxDO[21]) );
  XOR2_X1 output_mapping_2_U5 ( .A(InvUnmappedxD[19]), .B(InvUnmappedxD[21]), 
        .Z(QxDO[23]) );
  XNOR2_X1 output_mapping_2_U4 ( .A(output_mapping_2_n7), .B(InvUnmappedxD[17]), .ZN(QxDO[17]) );
  XNOR2_X1 output_mapping_2_U3 ( .A(InvUnmappedxD[21]), .B(InvUnmappedxD[20]), 
        .ZN(output_mapping_2_n7) );
  XNOR2_X1 output_mapping_2_U2 ( .A(InvUnmappedxD[17]), .B(output_mapping_2_n9), .ZN(QxDO[16]) );
  XNOR2_X1 output_mapping_2_U1 ( .A(InvUnmappedxD[22]), .B(InvUnmappedxD[20]), 
        .ZN(output_mapping_2_n9) );
  XNOR2_X1 input_mapping_1_U14 ( .A(input_mapping_1_n23), .B(
        input_mapping_1_n22), .ZN(mappedxD_1__7_) );
  XOR2_X1 input_mapping_1_U13 ( .A(XxDI[12]), .B(mappedxD_1__1_), .Z(
        mappedxD_1__6_) );
  XNOR2_X1 input_mapping_1_U12 ( .A(input_mapping_1_n21), .B(
        input_mapping_1_n20), .ZN(mappedxD_1__5_) );
  XNOR2_X1 input_mapping_1_U11 ( .A(XxDI[8]), .B(input_mapping_1_n22), .ZN(
        mappedxD_1__4_) );
  XNOR2_X1 input_mapping_1_U10 ( .A(XxDI[15]), .B(input_mapping_1_n21), .ZN(
        input_mapping_1_n22) );
  XNOR2_X1 input_mapping_1_U9 ( .A(input_mapping_1_n19), .B(
        input_mapping_1_n18), .ZN(mappedxD_1__3_) );
  XNOR2_X1 input_mapping_1_U8 ( .A(input_mapping_1_n20), .B(XxDI[11]), .ZN(
        input_mapping_1_n18) );
  XNOR2_X1 input_mapping_1_U7 ( .A(XxDI[15]), .B(XxDI[12]), .ZN(
        input_mapping_1_n19) );
  XOR2_X1 input_mapping_1_U6 ( .A(XxDI[8]), .B(input_mapping_1_n21), .Z(
        mappedxD_1__1_) );
  XOR2_X1 input_mapping_1_U5 ( .A(XxDI[14]), .B(XxDI[13]), .Z(
        input_mapping_1_n21) );
  XNOR2_X1 input_mapping_1_U4 ( .A(input_mapping_1_n23), .B(
        input_mapping_1_n17), .ZN(mappedxD_1__0_) );
  XNOR2_X1 input_mapping_1_U3 ( .A(XxDI[14]), .B(XxDI[11]), .ZN(
        input_mapping_1_n17) );
  XNOR2_X1 input_mapping_1_U2 ( .A(XxDI[10]), .B(input_mapping_1_n20), .ZN(
        input_mapping_1_n23) );
  XNOR2_X1 input_mapping_1_U1 ( .A(XxDI[8]), .B(XxDI[9]), .ZN(
        input_mapping_1_n20) );
  XOR2_X1 square_scaler_gf24_1_U3 ( .A(Y0xorY12xD[4]), .B(Y0xorY1xD[4]), .Z(
        Y0xorY12xD[7]) );
  XOR2_X1 square_scaler_gf24_1_U2 ( .A(Y0xorY1xD[3]), .B(Y0xorY1xD[5]), .Z(
        Y0xorY12xD[6]) );
  XOR2_X1 square_scaler_gf24_1_U1 ( .A(Y0xorY12xD[4]), .B(Y0xorY1xD[3]), .Z(
        Y0xorY12xD[5]) );
  XOR2_X1 output_mapping_1_U11 ( .A(InvUnmappedxD[11]), .B(InvUnmappedxD[15]), 
        .Z(QxDO[14]) );
  XNOR2_X1 output_mapping_1_U10 ( .A(QxDO[12]), .B(output_mapping_1_n9), .ZN(
        QxDO[11]) );
  XOR2_X1 output_mapping_1_U9 ( .A(QxDO[15]), .B(InvUnmappedxD[15]), .Z(
        QxDO[12]) );
  XNOR2_X1 output_mapping_1_U8 ( .A(output_mapping_1_n8), .B(QxDO[13]), .ZN(
        QxDO[10]) );
  XNOR2_X1 output_mapping_1_U7 ( .A(QxDO[15]), .B(InvUnmappedxD[10]), .ZN(
        output_mapping_1_n8) );
  XOR2_X1 output_mapping_1_U6 ( .A(InvUnmappedxD[14]), .B(InvUnmappedxD[8]), 
        .Z(QxDO[13]) );
  XOR2_X1 output_mapping_1_U5 ( .A(InvUnmappedxD[11]), .B(InvUnmappedxD[13]), 
        .Z(QxDO[15]) );
  XNOR2_X1 output_mapping_1_U4 ( .A(output_mapping_1_n7), .B(InvUnmappedxD[9]), 
        .ZN(QxDO[9]) );
  XNOR2_X1 output_mapping_1_U3 ( .A(InvUnmappedxD[13]), .B(InvUnmappedxD[12]), 
        .ZN(output_mapping_1_n7) );
  XNOR2_X1 output_mapping_1_U2 ( .A(InvUnmappedxD[9]), .B(output_mapping_1_n9), 
        .ZN(QxDO[8]) );
  XNOR2_X1 output_mapping_1_U1 ( .A(InvUnmappedxD[14]), .B(InvUnmappedxD[12]), 
        .ZN(output_mapping_1_n9) );
  XNOR2_X1 input_mapping_0_U14 ( .A(input_mapping_0_n23), .B(
        input_mapping_0_n22), .ZN(mappedxD_0__7_) );
  XOR2_X1 input_mapping_0_U13 ( .A(XxDI[4]), .B(mappedxD_0__1_), .Z(
        mappedxD_0__6_) );
  XNOR2_X1 input_mapping_0_U12 ( .A(input_mapping_0_n21), .B(
        input_mapping_0_n20), .ZN(mappedxD_0__5_) );
  XNOR2_X1 input_mapping_0_U11 ( .A(XxDI[0]), .B(input_mapping_0_n22), .ZN(
        mappedxD_0__4_) );
  XNOR2_X1 input_mapping_0_U10 ( .A(XxDI[7]), .B(input_mapping_0_n21), .ZN(
        input_mapping_0_n22) );
  XNOR2_X1 input_mapping_0_U9 ( .A(input_mapping_0_n19), .B(
        input_mapping_0_n18), .ZN(mappedxD_0__3_) );
  XNOR2_X1 input_mapping_0_U8 ( .A(input_mapping_0_n20), .B(XxDI[3]), .ZN(
        input_mapping_0_n18) );
  XNOR2_X1 input_mapping_0_U7 ( .A(XxDI[7]), .B(XxDI[4]), .ZN(
        input_mapping_0_n19) );
  XOR2_X1 input_mapping_0_U6 ( .A(XxDI[0]), .B(input_mapping_0_n21), .Z(
        mappedxD_0__1_) );
  XOR2_X1 input_mapping_0_U5 ( .A(XxDI[6]), .B(XxDI[5]), .Z(
        input_mapping_0_n21) );
  XNOR2_X1 input_mapping_0_U4 ( .A(input_mapping_0_n23), .B(
        input_mapping_0_n17), .ZN(mappedxD_0__0_) );
  XNOR2_X1 input_mapping_0_U3 ( .A(XxDI[6]), .B(XxDI[3]), .ZN(
        input_mapping_0_n17) );
  XNOR2_X1 input_mapping_0_U2 ( .A(XxDI[2]), .B(input_mapping_0_n20), .ZN(
        input_mapping_0_n23) );
  XNOR2_X1 input_mapping_0_U1 ( .A(XxDI[0]), .B(XxDI[1]), .ZN(
        input_mapping_0_n20) );
  XOR2_X1 square_scaler_gf24_0_U3 ( .A(Y0xorY12xD[0]), .B(Y0xorY1xD[1]), .Z(
        Y0xorY12xD[3]) );
  XOR2_X1 square_scaler_gf24_0_U2 ( .A(Y0xorY1xD[0]), .B(Y0xorY1xD[2]), .Z(
        Y0xorY12xD[2]) );
  XOR2_X1 square_scaler_gf24_0_U1 ( .A(Y0xorY12xD[0]), .B(Y0xorY1xD[0]), .Z(
        Y0xorY12xD[1]) );
  XOR2_X1 output_mapping_0_U11 ( .A(InvUnmappedxD[3]), .B(InvUnmappedxD[7]), 
        .Z(InvMappedxD_0__6_) );
  XNOR2_X1 output_mapping_0_U10 ( .A(QxDO[4]), .B(output_mapping_0_n9), .ZN(
        QxDO[3]) );
  XOR2_X1 output_mapping_0_U9 ( .A(QxDO[7]), .B(InvUnmappedxD[7]), .Z(QxDO[4])
         );
  XNOR2_X1 output_mapping_0_U8 ( .A(output_mapping_0_n8), .B(InvMappedxD_0__5_), .ZN(QxDO[2]) );
  XNOR2_X1 output_mapping_0_U7 ( .A(QxDO[7]), .B(InvUnmappedxD[2]), .ZN(
        output_mapping_0_n8) );
  XOR2_X1 output_mapping_0_U6 ( .A(InvUnmappedxD[6]), .B(InvUnmappedxD[0]), 
        .Z(InvMappedxD_0__5_) );
  XOR2_X1 output_mapping_0_U5 ( .A(InvUnmappedxD[3]), .B(InvUnmappedxD[5]), 
        .Z(QxDO[7]) );
  XNOR2_X1 output_mapping_0_U4 ( .A(output_mapping_0_n7), .B(InvUnmappedxD[1]), 
        .ZN(InvMappedxD_0__1_) );
  XNOR2_X1 output_mapping_0_U3 ( .A(InvUnmappedxD[5]), .B(InvUnmappedxD[4]), 
        .ZN(output_mapping_0_n7) );
  XNOR2_X1 output_mapping_0_U2 ( .A(InvUnmappedxD[1]), .B(output_mapping_0_n9), 
        .ZN(InvMappedxD_0__0_) );
  XNOR2_X1 output_mapping_0_U1 ( .A(InvUnmappedxD[6]), .B(InvUnmappedxD[4]), 
        .ZN(output_mapping_0_n9) );
  XNOR2_X1 mul_y0y1_U98 ( .A(mul_y0y1_n32), .B(mul_y0y1_n31), .ZN(
        Y0mulY1xD[15]) );
  XNOR2_X1 mul_y0y1_U97 ( .A(mul_y0y1_n34), .B(mul_y0y1_n33), .ZN(mul_y0y1_n31) );
  XOR2_X1 mul_y0y1_U96 ( .A(mul_y0y1_n36), .B(mul_y0y1_n35), .Z(mul_y0y1_n32)
         );
  XNOR2_X1 mul_y0y1_U95 ( .A(mul_y0y1_n30), .B(mul_y0y1_n29), .ZN(
        Y0mulY1xD[14]) );
  XNOR2_X1 mul_y0y1_U94 ( .A(mul_y0y1_n38), .B(mul_y0y1_n37), .ZN(mul_y0y1_n29) );
  XOR2_X1 mul_y0y1_U93 ( .A(mul_y0y1_n40), .B(mul_y0y1_n39), .Z(mul_y0y1_n30)
         );
  XNOR2_X1 mul_y0y1_U92 ( .A(mul_y0y1_n28), .B(mul_y0y1_n27), .ZN(
        Y0mulY1xD[13]) );
  XNOR2_X1 mul_y0y1_U91 ( .A(mul_y0y1_n42), .B(mul_y0y1_n41), .ZN(mul_y0y1_n27) );
  XOR2_X1 mul_y0y1_U90 ( .A(mul_y0y1_n44), .B(mul_y0y1_n43), .Z(mul_y0y1_n28)
         );
  XNOR2_X1 mul_y0y1_U89 ( .A(mul_y0y1_n26), .B(mul_y0y1_n25), .ZN(
        Y0mulY1xD[12]) );
  XNOR2_X1 mul_y0y1_U88 ( .A(mul_y0y1_n46), .B(mul_y0y1_n45), .ZN(mul_y0y1_n25) );
  XOR2_X1 mul_y0y1_U87 ( .A(mul_y0y1_n48), .B(mul_y0y1_n47), .Z(mul_y0y1_n26)
         );
  XNOR2_X1 mul_y0y1_U86 ( .A(mul_y0y1_n24), .B(mul_y0y1_n23), .ZN(
        Y0mulY1xD[11]) );
  XNOR2_X1 mul_y0y1_U85 ( .A(mul_y0y1_n50), .B(mul_y0y1_n49), .ZN(mul_y0y1_n23) );
  XOR2_X1 mul_y0y1_U84 ( .A(mul_y0y1_n52), .B(mul_y0y1_n51), .Z(mul_y0y1_n24)
         );
  XNOR2_X1 mul_y0y1_U83 ( .A(mul_y0y1_n22), .B(mul_y0y1_n21), .ZN(
        Y0mulY1xD[10]) );
  XNOR2_X1 mul_y0y1_U82 ( .A(mul_y0y1_n54), .B(mul_y0y1_n53), .ZN(mul_y0y1_n21) );
  XOR2_X1 mul_y0y1_U81 ( .A(mul_y0y1_n56), .B(mul_y0y1_n55), .Z(mul_y0y1_n22)
         );
  XNOR2_X1 mul_y0y1_U80 ( .A(mul_y0y1_n20), .B(mul_y0y1_n19), .ZN(Y0mulY1xD[9]) );
  XNOR2_X1 mul_y0y1_U79 ( .A(mul_y0y1_n58), .B(mul_y0y1_n57), .ZN(mul_y0y1_n19) );
  XOR2_X1 mul_y0y1_U78 ( .A(mul_y0y1_n60), .B(mul_y0y1_n59), .Z(mul_y0y1_n20)
         );
  XNOR2_X1 mul_y0y1_U77 ( .A(mul_y0y1_n18), .B(mul_y0y1_n17), .ZN(Y0mulY1xD[8]) );
  XNOR2_X1 mul_y0y1_U76 ( .A(mul_y0y1_n62), .B(mul_y0y1_n61), .ZN(mul_y0y1_n17) );
  XOR2_X1 mul_y0y1_U75 ( .A(mul_y0y1_n64), .B(mul_y0y1_n63), .Z(mul_y0y1_n18)
         );
  XNOR2_X1 mul_y0y1_U74 ( .A(mul_y0y1_n16), .B(mul_y0y1_n15), .ZN(Y0mulY1xD[7]) );
  XNOR2_X1 mul_y0y1_U73 ( .A(mul_y0y1_n66), .B(mul_y0y1_n65), .ZN(mul_y0y1_n15) );
  XOR2_X1 mul_y0y1_U72 ( .A(mul_y0y1_n68), .B(mul_y0y1_n67), .Z(mul_y0y1_n16)
         );
  XNOR2_X1 mul_y0y1_U71 ( .A(mul_y0y1_n14), .B(mul_y0y1_n13), .ZN(Y0mulY1xD[6]) );
  XNOR2_X1 mul_y0y1_U70 ( .A(mul_y0y1_n70), .B(mul_y0y1_n69), .ZN(mul_y0y1_n13) );
  XOR2_X1 mul_y0y1_U69 ( .A(mul_y0y1_n72), .B(mul_y0y1_n71), .Z(mul_y0y1_n14)
         );
  XNOR2_X1 mul_y0y1_U68 ( .A(mul_y0y1_n12), .B(mul_y0y1_n11), .ZN(Y0mulY1xD[5]) );
  XNOR2_X1 mul_y0y1_U67 ( .A(mul_y0y1_n74), .B(mul_y0y1_n73), .ZN(mul_y0y1_n11) );
  XOR2_X1 mul_y0y1_U66 ( .A(mul_y0y1_n76), .B(mul_y0y1_n75), .Z(mul_y0y1_n12)
         );
  XNOR2_X1 mul_y0y1_U65 ( .A(mul_y0y1_n10), .B(mul_y0y1_n9), .ZN(Y0mulY1xD[4])
         );
  XNOR2_X1 mul_y0y1_U64 ( .A(mul_y0y1_n78), .B(mul_y0y1_n77), .ZN(mul_y0y1_n9)
         );
  XOR2_X1 mul_y0y1_U63 ( .A(mul_y0y1_n80), .B(mul_y0y1_n79), .Z(mul_y0y1_n10)
         );
  XNOR2_X1 mul_y0y1_U62 ( .A(mul_y0y1_n8), .B(mul_y0y1_n7), .ZN(Y0mulY1xD[3])
         );
  XNOR2_X1 mul_y0y1_U61 ( .A(mul_y0y1_n82), .B(mul_y0y1_n81), .ZN(mul_y0y1_n7)
         );
  XOR2_X1 mul_y0y1_U60 ( .A(mul_y0y1_n84), .B(mul_y0y1_n83), .Z(mul_y0y1_n8)
         );
  XNOR2_X1 mul_y0y1_U59 ( .A(mul_y0y1_n6), .B(mul_y0y1_n5), .ZN(Y0mulY1xD[2])
         );
  XNOR2_X1 mul_y0y1_U58 ( .A(mul_y0y1_n86), .B(mul_y0y1_n85), .ZN(mul_y0y1_n5)
         );
  XOR2_X1 mul_y0y1_U57 ( .A(mul_y0y1_n88), .B(mul_y0y1_n87), .Z(mul_y0y1_n6)
         );
  XNOR2_X1 mul_y0y1_U56 ( .A(mul_y0y1_n4), .B(mul_y0y1_n3), .ZN(Y0mulY1xD[1])
         );
  XNOR2_X1 mul_y0y1_U55 ( .A(mul_y0y1_n90), .B(mul_y0y1_n89), .ZN(mul_y0y1_n3)
         );
  XOR2_X1 mul_y0y1_U54 ( .A(mul_y0y1_n92), .B(mul_y0y1_n91), .Z(mul_y0y1_n4)
         );
  XNOR2_X1 mul_y0y1_U53 ( .A(mul_y0y1_n2), .B(mul_y0y1_n1), .ZN(Y0mulY1xD[0])
         );
  XNOR2_X1 mul_y0y1_U52 ( .A(mul_y0y1_n94), .B(mul_y0y1_n93), .ZN(mul_y0y1_n1)
         );
  XOR2_X1 mul_y0y1_U51 ( .A(mul_y0y1_n96), .B(mul_y0y1_n95), .Z(mul_y0y1_n2)
         );
  XOR2_X1 mul_y0y1_U50 ( .A(Zmul1xDI[11]), .B(mul_y0y1_Xi_mul_Yj_9__3_), .Z(
        mul_y0y1_FFxDN[39]) );
  XOR2_X1 mul_y0y1_U49 ( .A(Zmul1xDI[10]), .B(mul_y0y1_Xi_mul_Yj_9__2_), .Z(
        mul_y0y1_FFxDN[38]) );
  XOR2_X1 mul_y0y1_U48 ( .A(Zmul1xDI[9]), .B(mul_y0y1_Xi_mul_Yj_9__1_), .Z(
        mul_y0y1_FFxDN[37]) );
  XOR2_X1 mul_y0y1_U47 ( .A(Zmul1xDI[8]), .B(mul_y0y1_Xi_mul_Yj_9__0_), .Z(
        mul_y0y1_FFxDN[36]) );
  XOR2_X1 mul_y0y1_U46 ( .A(Zmul1xDI[7]), .B(mul_y0y1_Xi_mul_Yj_8__3_), .Z(
        mul_y0y1_FFxDN[35]) );
  XOR2_X1 mul_y0y1_U45 ( .A(Zmul1xDI[6]), .B(mul_y0y1_Xi_mul_Yj_8__2_), .Z(
        mul_y0y1_FFxDN[34]) );
  XOR2_X1 mul_y0y1_U44 ( .A(Zmul1xDI[5]), .B(mul_y0y1_Xi_mul_Yj_8__1_), .Z(
        mul_y0y1_FFxDN[33]) );
  XOR2_X1 mul_y0y1_U43 ( .A(Zmul1xDI[4]), .B(mul_y0y1_Xi_mul_Yj_8__0_), .Z(
        mul_y0y1_FFxDN[32]) );
  XOR2_X1 mul_y0y1_U42 ( .A(Zmul1xDI[19]), .B(mul_y0y1_Xi_mul_Yj_7__3_), .Z(
        mul_y0y1_FFxDN[31]) );
  XOR2_X1 mul_y0y1_U41 ( .A(Zmul1xDI[18]), .B(mul_y0y1_Xi_mul_Yj_7__2_), .Z(
        mul_y0y1_FFxDN[30]) );
  XOR2_X1 mul_y0y1_U40 ( .A(Zmul1xDI[17]), .B(mul_y0y1_Xi_mul_Yj_7__1_), .Z(
        mul_y0y1_FFxDN[29]) );
  XOR2_X1 mul_y0y1_U39 ( .A(Zmul1xDI[16]), .B(mul_y0y1_Xi_mul_Yj_7__0_), .Z(
        mul_y0y1_FFxDN[28]) );
  XOR2_X1 mul_y0y1_U38 ( .A(Zmul1xDI[11]), .B(mul_y0y1_Xi_mul_Yj_6__3_), .Z(
        mul_y0y1_FFxDN[27]) );
  XOR2_X1 mul_y0y1_U37 ( .A(Zmul1xDI[10]), .B(mul_y0y1_Xi_mul_Yj_6__2_), .Z(
        mul_y0y1_FFxDN[26]) );
  XOR2_X1 mul_y0y1_U36 ( .A(Zmul1xDI[9]), .B(mul_y0y1_Xi_mul_Yj_6__1_), .Z(
        mul_y0y1_FFxDN[25]) );
  XOR2_X1 mul_y0y1_U35 ( .A(Zmul1xDI[8]), .B(mul_y0y1_Xi_mul_Yj_6__0_), .Z(
        mul_y0y1_FFxDN[24]) );
  XOR2_X1 mul_y0y1_U34 ( .A(Zmul1xDI[3]), .B(mul_y0y1_Xi_mul_Yj_4__3_), .Z(
        mul_y0y1_FFxDN[19]) );
  XOR2_X1 mul_y0y1_U33 ( .A(Zmul1xDI[2]), .B(mul_y0y1_Xi_mul_Yj_4__2_), .Z(
        mul_y0y1_FFxDN[18]) );
  XOR2_X1 mul_y0y1_U32 ( .A(Zmul1xDI[1]), .B(mul_y0y1_Xi_mul_Yj_4__1_), .Z(
        mul_y0y1_FFxDN[17]) );
  XOR2_X1 mul_y0y1_U31 ( .A(Zmul1xDI[0]), .B(mul_y0y1_Xi_mul_Yj_4__0_), .Z(
        mul_y0y1_FFxDN[16]) );
  XOR2_X1 mul_y0y1_U30 ( .A(Zmul1xDI[15]), .B(mul_y0y1_Xi_mul_Yj_3__3_), .Z(
        mul_y0y1_FFxDN[15]) );
  XOR2_X1 mul_y0y1_U29 ( .A(Zmul1xDI[14]), .B(mul_y0y1_Xi_mul_Yj_3__2_), .Z(
        mul_y0y1_FFxDN[14]) );
  XOR2_X1 mul_y0y1_U28 ( .A(Zmul1xDI[13]), .B(mul_y0y1_Xi_mul_Yj_3__1_), .Z(
        mul_y0y1_FFxDN[13]) );
  XOR2_X1 mul_y0y1_U27 ( .A(Zmul1xDI[12]), .B(mul_y0y1_Xi_mul_Yj_3__0_), .Z(
        mul_y0y1_FFxDN[12]) );
  XOR2_X1 mul_y0y1_U26 ( .A(Zmul1xDI[7]), .B(mul_y0y1_Xi_mul_Yj_2__3_), .Z(
        mul_y0y1_FFxDN[11]) );
  XOR2_X1 mul_y0y1_U25 ( .A(Zmul1xDI[6]), .B(mul_y0y1_Xi_mul_Yj_2__2_), .Z(
        mul_y0y1_FFxDN[10]) );
  XOR2_X1 mul_y0y1_U24 ( .A(Zmul1xDI[5]), .B(mul_y0y1_Xi_mul_Yj_2__1_), .Z(
        mul_y0y1_FFxDN[9]) );
  XOR2_X1 mul_y0y1_U23 ( .A(Zmul1xDI[4]), .B(mul_y0y1_Xi_mul_Yj_2__0_), .Z(
        mul_y0y1_FFxDN[8]) );
  XOR2_X1 mul_y0y1_U22 ( .A(Zmul1xDI[3]), .B(mul_y0y1_Xi_mul_Yj_1__3_), .Z(
        mul_y0y1_FFxDN[7]) );
  XOR2_X1 mul_y0y1_U21 ( .A(Zmul1xDI[2]), .B(mul_y0y1_Xi_mul_Yj_1__2_), .Z(
        mul_y0y1_FFxDN[6]) );
  XOR2_X1 mul_y0y1_U20 ( .A(Zmul1xDI[1]), .B(mul_y0y1_Xi_mul_Yj_1__1_), .Z(
        mul_y0y1_FFxDN[5]) );
  XOR2_X1 mul_y0y1_U19 ( .A(Zmul1xDI[0]), .B(mul_y0y1_Xi_mul_Yj_1__0_), .Z(
        mul_y0y1_FFxDN[4]) );
  XOR2_X1 mul_y0y1_U18 ( .A(Zmul1xDI[23]), .B(mul_y0y1_Xi_mul_Yj_14__3_), .Z(
        mul_y0y1_FFxDN[59]) );
  XOR2_X1 mul_y0y1_U17 ( .A(Zmul1xDI[22]), .B(mul_y0y1_Xi_mul_Yj_14__2_), .Z(
        mul_y0y1_FFxDN[58]) );
  XOR2_X1 mul_y0y1_U16 ( .A(Zmul1xDI[21]), .B(mul_y0y1_Xi_mul_Yj_14__1_), .Z(
        mul_y0y1_FFxDN[57]) );
  XOR2_X1 mul_y0y1_U15 ( .A(Zmul1xDI[20]), .B(mul_y0y1_Xi_mul_Yj_14__0_), .Z(
        mul_y0y1_FFxDN[56]) );
  XOR2_X1 mul_y0y1_U14 ( .A(Zmul1xDI[19]), .B(mul_y0y1_Xi_mul_Yj_13__3_), .Z(
        mul_y0y1_FFxDN[55]) );
  XOR2_X1 mul_y0y1_U13 ( .A(Zmul1xDI[18]), .B(mul_y0y1_Xi_mul_Yj_13__2_), .Z(
        mul_y0y1_FFxDN[54]) );
  XOR2_X1 mul_y0y1_U12 ( .A(Zmul1xDI[17]), .B(mul_y0y1_Xi_mul_Yj_13__1_), .Z(
        mul_y0y1_FFxDN[53]) );
  XOR2_X1 mul_y0y1_U11 ( .A(Zmul1xDI[16]), .B(mul_y0y1_Xi_mul_Yj_13__0_), .Z(
        mul_y0y1_FFxDN[52]) );
  XOR2_X1 mul_y0y1_U10 ( .A(Zmul1xDI[15]), .B(mul_y0y1_Xi_mul_Yj_12__3_), .Z(
        mul_y0y1_FFxDN[51]) );
  XOR2_X1 mul_y0y1_U9 ( .A(Zmul1xDI[14]), .B(mul_y0y1_Xi_mul_Yj_12__2_), .Z(
        mul_y0y1_FFxDN[50]) );
  XOR2_X1 mul_y0y1_U8 ( .A(Zmul1xDI[13]), .B(mul_y0y1_Xi_mul_Yj_12__1_), .Z(
        mul_y0y1_FFxDN[49]) );
  XOR2_X1 mul_y0y1_U7 ( .A(Zmul1xDI[12]), .B(mul_y0y1_Xi_mul_Yj_12__0_), .Z(
        mul_y0y1_FFxDN[48]) );
  XOR2_X1 mul_y0y1_U6 ( .A(Zmul1xDI[23]), .B(mul_y0y1_Xi_mul_Yj_11__3_), .Z(
        mul_y0y1_FFxDN[47]) );
  XOR2_X1 mul_y0y1_U5 ( .A(Zmul1xDI[22]), .B(mul_y0y1_Xi_mul_Yj_11__2_), .Z(
        mul_y0y1_FFxDN[46]) );
  XOR2_X1 mul_y0y1_U4 ( .A(Zmul1xDI[21]), .B(mul_y0y1_Xi_mul_Yj_11__1_), .Z(
        mul_y0y1_FFxDN[45]) );
  XOR2_X1 mul_y0y1_U3 ( .A(Zmul1xDI[20]), .B(mul_y0y1_Xi_mul_Yj_11__0_), .Z(
        mul_y0y1_FFxDN[44]) );
  DFF_X1 mul_y0y1_FFxDP_reg_1__3_ ( .D(mul_y0y1_FFxDN[7]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n84) );
  DFF_X1 mul_y0y1_FFxDP_reg_2__3_ ( .D(mul_y0y1_FFxDN[11]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n81) );
  DFF_X1 mul_y0y1_FFxDP_reg_3__3_ ( .D(mul_y0y1_FFxDN[15]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n82) );
  DFF_X1 mul_y0y1_FFxDP_reg_4__3_ ( .D(mul_y0y1_FFxDN[19]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n67) );
  DFF_X1 mul_y0y1_FFxDP_reg_6__3_ ( .D(mul_y0y1_FFxDN[27]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n65) );
  DFF_X1 mul_y0y1_FFxDP_reg_7__3_ ( .D(mul_y0y1_FFxDN[31]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n66) );
  DFF_X1 mul_y0y1_FFxDP_reg_8__3_ ( .D(mul_y0y1_FFxDN[35]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n49) );
  DFF_X1 mul_y0y1_FFxDP_reg_9__3_ ( .D(mul_y0y1_FFxDN[39]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n50) );
  DFF_X1 mul_y0y1_FFxDP_reg_11__3_ ( .D(mul_y0y1_FFxDN[47]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n52) );
  DFF_X1 mul_y0y1_FFxDP_reg_12__3_ ( .D(mul_y0y1_FFxDN[51]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n35) );
  DFF_X1 mul_y0y1_FFxDP_reg_13__3_ ( .D(mul_y0y1_FFxDN[55]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n36) );
  DFF_X1 mul_y0y1_FFxDP_reg_14__3_ ( .D(mul_y0y1_FFxDN[59]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n33) );
  DFF_X1 mul_y0y1_FFxDP_reg_1__1_ ( .D(mul_y0y1_FFxDN[5]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n92) );
  DFF_X1 mul_y0y1_FFxDP_reg_2__1_ ( .D(mul_y0y1_FFxDN[9]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n89) );
  DFF_X1 mul_y0y1_FFxDP_reg_3__1_ ( .D(mul_y0y1_FFxDN[13]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n90) );
  DFF_X1 mul_y0y1_FFxDP_reg_4__1_ ( .D(mul_y0y1_FFxDN[17]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n75) );
  DFF_X1 mul_y0y1_FFxDP_reg_6__1_ ( .D(mul_y0y1_FFxDN[25]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n73) );
  DFF_X1 mul_y0y1_FFxDP_reg_7__1_ ( .D(mul_y0y1_FFxDN[29]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n74) );
  DFF_X1 mul_y0y1_FFxDP_reg_8__1_ ( .D(mul_y0y1_FFxDN[33]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n57) );
  DFF_X1 mul_y0y1_FFxDP_reg_9__1_ ( .D(mul_y0y1_FFxDN[37]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n58) );
  DFF_X1 mul_y0y1_FFxDP_reg_11__1_ ( .D(mul_y0y1_FFxDN[45]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n60) );
  DFF_X1 mul_y0y1_FFxDP_reg_12__1_ ( .D(mul_y0y1_FFxDN[49]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n43) );
  DFF_X1 mul_y0y1_FFxDP_reg_13__1_ ( .D(mul_y0y1_FFxDN[53]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n44) );
  DFF_X1 mul_y0y1_FFxDP_reg_14__1_ ( .D(mul_y0y1_FFxDN[57]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n41) );
  DFF_X1 mul_y0y1_FFxDP_reg_1__2_ ( .D(mul_y0y1_FFxDN[6]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n88) );
  DFF_X1 mul_y0y1_FFxDP_reg_2__2_ ( .D(mul_y0y1_FFxDN[10]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n85) );
  DFF_X1 mul_y0y1_FFxDP_reg_3__2_ ( .D(mul_y0y1_FFxDN[14]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n86) );
  DFF_X1 mul_y0y1_FFxDP_reg_4__2_ ( .D(mul_y0y1_FFxDN[18]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n71) );
  DFF_X1 mul_y0y1_FFxDP_reg_6__2_ ( .D(mul_y0y1_FFxDN[26]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n69) );
  DFF_X1 mul_y0y1_FFxDP_reg_7__2_ ( .D(mul_y0y1_FFxDN[30]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n70) );
  DFF_X1 mul_y0y1_FFxDP_reg_8__2_ ( .D(mul_y0y1_FFxDN[34]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n53) );
  DFF_X1 mul_y0y1_FFxDP_reg_9__2_ ( .D(mul_y0y1_FFxDN[38]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n54) );
  DFF_X1 mul_y0y1_FFxDP_reg_11__2_ ( .D(mul_y0y1_FFxDN[46]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n56) );
  DFF_X1 mul_y0y1_FFxDP_reg_12__2_ ( .D(mul_y0y1_FFxDN[50]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n39) );
  DFF_X1 mul_y0y1_FFxDP_reg_13__2_ ( .D(mul_y0y1_FFxDN[54]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n40) );
  DFF_X1 mul_y0y1_FFxDP_reg_14__2_ ( .D(mul_y0y1_FFxDN[58]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n37) );
  DFF_X1 mul_y0y1_FFxDP_reg_1__0_ ( .D(mul_y0y1_FFxDN[4]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n96) );
  DFF_X1 mul_y0y1_FFxDP_reg_2__0_ ( .D(mul_y0y1_FFxDN[8]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n93) );
  DFF_X1 mul_y0y1_FFxDP_reg_3__0_ ( .D(mul_y0y1_FFxDN[12]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n94) );
  DFF_X1 mul_y0y1_FFxDP_reg_4__0_ ( .D(mul_y0y1_FFxDN[16]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n79) );
  DFF_X1 mul_y0y1_FFxDP_reg_6__0_ ( .D(mul_y0y1_FFxDN[24]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n77) );
  DFF_X1 mul_y0y1_FFxDP_reg_7__0_ ( .D(mul_y0y1_FFxDN[28]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n78) );
  DFF_X1 mul_y0y1_FFxDP_reg_8__0_ ( .D(mul_y0y1_FFxDN[32]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n61) );
  DFF_X1 mul_y0y1_FFxDP_reg_9__0_ ( .D(mul_y0y1_FFxDN[36]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n62) );
  DFF_X1 mul_y0y1_FFxDP_reg_11__0_ ( .D(mul_y0y1_FFxDN[44]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n64) );
  DFF_X1 mul_y0y1_FFxDP_reg_12__0_ ( .D(mul_y0y1_FFxDN[48]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n47) );
  DFF_X1 mul_y0y1_FFxDP_reg_13__0_ ( .D(mul_y0y1_FFxDN[52]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n48) );
  DFF_X1 mul_y0y1_FFxDP_reg_14__0_ ( .D(mul_y0y1_FFxDN[56]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n45) );
  DFF_X1 mul_y0y1_FFxDP_reg_0__3_ ( .D(mul_y0y1_FFxDN[3]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n83) );
  DFF_X1 mul_y0y1_FFxDP_reg_5__3_ ( .D(mul_y0y1_FFxDN[23]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n68) );
  DFF_X1 mul_y0y1_FFxDP_reg_10__3_ ( .D(mul_y0y1_FFxDN[43]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n51) );
  DFF_X1 mul_y0y1_FFxDP_reg_15__3_ ( .D(mul_y0y1_FFxDN[63]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n34) );
  DFF_X1 mul_y0y1_FFxDP_reg_0__1_ ( .D(mul_y0y1_FFxDN[1]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n91) );
  DFF_X1 mul_y0y1_FFxDP_reg_5__1_ ( .D(mul_y0y1_FFxDN[21]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n76) );
  DFF_X1 mul_y0y1_FFxDP_reg_10__1_ ( .D(mul_y0y1_FFxDN[41]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n59) );
  DFF_X1 mul_y0y1_FFxDP_reg_15__1_ ( .D(mul_y0y1_FFxDN[61]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n42) );
  DFF_X1 mul_y0y1_FFxDP_reg_0__2_ ( .D(mul_y0y1_FFxDN[2]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n87) );
  DFF_X1 mul_y0y1_FFxDP_reg_5__2_ ( .D(mul_y0y1_FFxDN[22]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n72) );
  DFF_X1 mul_y0y1_FFxDP_reg_10__2_ ( .D(mul_y0y1_FFxDN[42]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n55) );
  DFF_X1 mul_y0y1_FFxDP_reg_15__2_ ( .D(mul_y0y1_FFxDN[62]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n38) );
  DFF_X1 mul_y0y1_FFxDP_reg_0__0_ ( .D(mul_y0y1_FFxDN[0]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n95) );
  DFF_X1 mul_y0y1_FFxDP_reg_5__0_ ( .D(mul_y0y1_FFxDN[20]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n80) );
  DFF_X1 mul_y0y1_FFxDP_reg_10__0_ ( .D(mul_y0y1_FFxDN[40]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n63) );
  DFF_X1 mul_y0y1_FFxDP_reg_15__0_ ( .D(mul_y0y1_FFxDN[60]), .CK(ClkxCI), .Q(), 
        .QN(mul_y0y1_n46) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_3_U29 ( .A(mul_y0y1_gf4_mul_3_3_n77), .B(
        mul_y0y1_gf4_mul_3_3_n76), .ZN(mul_y0y1_FFxDN[63]) );
  NAND2_X1 mul_y0y1_gf4_mul_3_3_U28 ( .A1(Y1xD[15]), .A2(Y0xD[15]), .ZN(
        mul_y0y1_gf4_mul_3_3_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_3_3_U27 ( .A(mul_y0y1_gf4_mul_3_3_n75), .B(
        mul_y0y1_gf4_mul_3_3_n74), .Z(mul_y0y1_gf4_mul_3_3_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_3_U26 ( .A(mul_y0y1_gf4_mul_3_3_n73), .B(
        mul_y0y1_gf4_mul_3_3_n72), .ZN(mul_y0y1_FFxDN[62]) );
  NAND2_X1 mul_y0y1_gf4_mul_3_3_U25 ( .A1(Y1xD[14]), .A2(Y0xD[14]), .ZN(
        mul_y0y1_gf4_mul_3_3_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_3_3_U24 ( .A(mul_y0y1_gf4_mul_3_3_n74), .B(
        mul_y0y1_gf4_mul_3_3_n71), .Z(mul_y0y1_gf4_mul_3_3_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_3_3_U23 ( .A1(mul_y0y1_gf4_mul_3_3_n70), .A2(
        mul_y0y1_gf4_mul_3_3_n69), .ZN(mul_y0y1_gf4_mul_3_3_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_3_U22 ( .A(Y1xD[14]), .B(Y1xD[15]), .ZN(
        mul_y0y1_gf4_mul_3_3_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_3_U21 ( .A(Y0xD[14]), .B(Y0xD[15]), .ZN(
        mul_y0y1_gf4_mul_3_3_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_3_U20 ( .A(mul_y0y1_gf4_mul_3_3_n68), .B(
        mul_y0y1_gf4_mul_3_3_n67), .ZN(mul_y0y1_FFxDN[61]) );
  NAND2_X1 mul_y0y1_gf4_mul_3_3_U19 ( .A1(Y1xD[13]), .A2(Y0xD[13]), .ZN(
        mul_y0y1_gf4_mul_3_3_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_3_3_U18 ( .A(mul_y0y1_gf4_mul_3_3_n75), .B(
        mul_y0y1_gf4_mul_3_3_n66), .Z(mul_y0y1_gf4_mul_3_3_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_3_U17 ( .A(mul_y0y1_gf4_mul_3_3_n65), .B(
        mul_y0y1_gf4_mul_3_3_n64), .ZN(mul_y0y1_gf4_mul_3_3_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_3_3_U16 ( .A1(mul_y0y1_gf4_mul_3_3_n63), .A2(
        mul_y0y1_gf4_mul_3_3_n62), .ZN(mul_y0y1_gf4_mul_3_3_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_3_U15 ( .A(mul_y0y1_gf4_mul_3_3_n61), .B(
        mul_y0y1_gf4_mul_3_3_n60), .ZN(mul_y0y1_gf4_mul_3_3_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_3_U14 ( .A(mul_y0y1_gf4_mul_3_3_n59), .B(
        mul_y0y1_gf4_mul_3_3_n58), .ZN(mul_y0y1_gf4_mul_3_3_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_3_U13 ( .A(mul_y0y1_gf4_mul_3_3_n57), .B(
        mul_y0y1_gf4_mul_3_3_n56), .ZN(mul_y0y1_FFxDN[60]) );
  NAND2_X1 mul_y0y1_gf4_mul_3_3_U12 ( .A1(Y1xD[12]), .A2(Y0xD[12]), .ZN(
        mul_y0y1_gf4_mul_3_3_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_3_3_U11 ( .A(mul_y0y1_gf4_mul_3_3_n66), .B(
        mul_y0y1_gf4_mul_3_3_n71), .Z(mul_y0y1_gf4_mul_3_3_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_3_U10 ( .A(mul_y0y1_gf4_mul_3_3_n55), .B(
        mul_y0y1_gf4_mul_3_3_n65), .ZN(mul_y0y1_gf4_mul_3_3_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_3_3_U9 ( .A1(mul_y0y1_gf4_mul_3_3_n61), .A2(
        mul_y0y1_gf4_mul_3_3_n59), .ZN(mul_y0y1_gf4_mul_3_3_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_3_U8 ( .A(Y1xD[12]), .B(Y1xD[14]), .ZN(
        mul_y0y1_gf4_mul_3_3_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_3_U7 ( .A(Y0xD[12]), .B(Y0xD[14]), .ZN(
        mul_y0y1_gf4_mul_3_3_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_3_3_U6 ( .A1(mul_y0y1_gf4_mul_3_3_n58), .A2(
        mul_y0y1_gf4_mul_3_3_n60), .ZN(mul_y0y1_gf4_mul_3_3_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_3_3_U5 ( .A(Y0xD[13]), .B(Y0xD[15]), .Z(
        mul_y0y1_gf4_mul_3_3_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_3_3_U4 ( .A(Y1xD[13]), .B(Y1xD[15]), .Z(
        mul_y0y1_gf4_mul_3_3_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_3_3_U3 ( .A1(mul_y0y1_gf4_mul_3_3_n54), .A2(
        mul_y0y1_gf4_mul_3_3_n53), .ZN(mul_y0y1_gf4_mul_3_3_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_3_U2 ( .A(Y1xD[12]), .B(Y1xD[13]), .ZN(
        mul_y0y1_gf4_mul_3_3_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_3_U1 ( .A(Y0xD[12]), .B(Y0xD[13]), .ZN(
        mul_y0y1_gf4_mul_3_3_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_2_U29 ( .A(mul_y0y1_gf4_mul_3_2_n77), .B(
        mul_y0y1_gf4_mul_3_2_n76), .ZN(mul_y0y1_Xi_mul_Yj_14__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_3_2_U28 ( .A1(Y1xD[15]), .A2(Y0xD[11]), .ZN(
        mul_y0y1_gf4_mul_3_2_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_3_2_U27 ( .A(mul_y0y1_gf4_mul_3_2_n75), .B(
        mul_y0y1_gf4_mul_3_2_n74), .Z(mul_y0y1_gf4_mul_3_2_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_2_U26 ( .A(mul_y0y1_gf4_mul_3_2_n73), .B(
        mul_y0y1_gf4_mul_3_2_n72), .ZN(mul_y0y1_Xi_mul_Yj_14__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_3_2_U25 ( .A1(Y1xD[14]), .A2(Y0xD[10]), .ZN(
        mul_y0y1_gf4_mul_3_2_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_3_2_U24 ( .A(mul_y0y1_gf4_mul_3_2_n74), .B(
        mul_y0y1_gf4_mul_3_2_n71), .Z(mul_y0y1_gf4_mul_3_2_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_3_2_U23 ( .A1(mul_y0y1_gf4_mul_3_2_n70), .A2(
        mul_y0y1_gf4_mul_3_2_n69), .ZN(mul_y0y1_gf4_mul_3_2_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_2_U22 ( .A(Y1xD[14]), .B(Y1xD[15]), .ZN(
        mul_y0y1_gf4_mul_3_2_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_2_U21 ( .A(Y0xD[10]), .B(Y0xD[11]), .ZN(
        mul_y0y1_gf4_mul_3_2_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_2_U20 ( .A(mul_y0y1_gf4_mul_3_2_n68), .B(
        mul_y0y1_gf4_mul_3_2_n67), .ZN(mul_y0y1_Xi_mul_Yj_14__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_3_2_U19 ( .A1(Y1xD[13]), .A2(Y0xD[9]), .ZN(
        mul_y0y1_gf4_mul_3_2_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_3_2_U18 ( .A(mul_y0y1_gf4_mul_3_2_n75), .B(
        mul_y0y1_gf4_mul_3_2_n66), .Z(mul_y0y1_gf4_mul_3_2_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_2_U17 ( .A(mul_y0y1_gf4_mul_3_2_n65), .B(
        mul_y0y1_gf4_mul_3_2_n64), .ZN(mul_y0y1_gf4_mul_3_2_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_3_2_U16 ( .A1(mul_y0y1_gf4_mul_3_2_n63), .A2(
        mul_y0y1_gf4_mul_3_2_n62), .ZN(mul_y0y1_gf4_mul_3_2_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_2_U15 ( .A(mul_y0y1_gf4_mul_3_2_n61), .B(
        mul_y0y1_gf4_mul_3_2_n60), .ZN(mul_y0y1_gf4_mul_3_2_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_2_U14 ( .A(mul_y0y1_gf4_mul_3_2_n59), .B(
        mul_y0y1_gf4_mul_3_2_n58), .ZN(mul_y0y1_gf4_mul_3_2_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_2_U13 ( .A(mul_y0y1_gf4_mul_3_2_n57), .B(
        mul_y0y1_gf4_mul_3_2_n56), .ZN(mul_y0y1_Xi_mul_Yj_14__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_3_2_U12 ( .A1(Y1xD[12]), .A2(Y0xD[8]), .ZN(
        mul_y0y1_gf4_mul_3_2_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_3_2_U11 ( .A(mul_y0y1_gf4_mul_3_2_n66), .B(
        mul_y0y1_gf4_mul_3_2_n71), .Z(mul_y0y1_gf4_mul_3_2_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_2_U10 ( .A(mul_y0y1_gf4_mul_3_2_n55), .B(
        mul_y0y1_gf4_mul_3_2_n65), .ZN(mul_y0y1_gf4_mul_3_2_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_3_2_U9 ( .A1(mul_y0y1_gf4_mul_3_2_n61), .A2(
        mul_y0y1_gf4_mul_3_2_n59), .ZN(mul_y0y1_gf4_mul_3_2_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_2_U8 ( .A(Y1xD[12]), .B(Y1xD[14]), .ZN(
        mul_y0y1_gf4_mul_3_2_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_2_U7 ( .A(Y0xD[8]), .B(Y0xD[10]), .ZN(
        mul_y0y1_gf4_mul_3_2_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_3_2_U6 ( .A1(mul_y0y1_gf4_mul_3_2_n58), .A2(
        mul_y0y1_gf4_mul_3_2_n60), .ZN(mul_y0y1_gf4_mul_3_2_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_3_2_U5 ( .A(Y0xD[9]), .B(Y0xD[11]), .Z(
        mul_y0y1_gf4_mul_3_2_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_3_2_U4 ( .A(Y1xD[13]), .B(Y1xD[15]), .Z(
        mul_y0y1_gf4_mul_3_2_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_3_2_U3 ( .A1(mul_y0y1_gf4_mul_3_2_n54), .A2(
        mul_y0y1_gf4_mul_3_2_n53), .ZN(mul_y0y1_gf4_mul_3_2_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_2_U2 ( .A(Y1xD[12]), .B(Y1xD[13]), .ZN(
        mul_y0y1_gf4_mul_3_2_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_2_U1 ( .A(Y0xD[8]), .B(Y0xD[9]), .ZN(
        mul_y0y1_gf4_mul_3_2_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_1_U29 ( .A(mul_y0y1_gf4_mul_3_1_n77), .B(
        mul_y0y1_gf4_mul_3_1_n76), .ZN(mul_y0y1_Xi_mul_Yj_13__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_3_1_U28 ( .A1(Y1xD[15]), .A2(Y0xD[7]), .ZN(
        mul_y0y1_gf4_mul_3_1_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_3_1_U27 ( .A(mul_y0y1_gf4_mul_3_1_n75), .B(
        mul_y0y1_gf4_mul_3_1_n74), .Z(mul_y0y1_gf4_mul_3_1_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_1_U26 ( .A(mul_y0y1_gf4_mul_3_1_n73), .B(
        mul_y0y1_gf4_mul_3_1_n72), .ZN(mul_y0y1_Xi_mul_Yj_13__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_3_1_U25 ( .A1(Y1xD[14]), .A2(Y0xD[6]), .ZN(
        mul_y0y1_gf4_mul_3_1_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_3_1_U24 ( .A(mul_y0y1_gf4_mul_3_1_n74), .B(
        mul_y0y1_gf4_mul_3_1_n71), .Z(mul_y0y1_gf4_mul_3_1_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_3_1_U23 ( .A1(mul_y0y1_gf4_mul_3_1_n70), .A2(
        mul_y0y1_gf4_mul_3_1_n69), .ZN(mul_y0y1_gf4_mul_3_1_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_1_U22 ( .A(Y1xD[14]), .B(Y1xD[15]), .ZN(
        mul_y0y1_gf4_mul_3_1_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_1_U21 ( .A(Y0xD[6]), .B(Y0xD[7]), .ZN(
        mul_y0y1_gf4_mul_3_1_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_1_U20 ( .A(mul_y0y1_gf4_mul_3_1_n68), .B(
        mul_y0y1_gf4_mul_3_1_n67), .ZN(mul_y0y1_Xi_mul_Yj_13__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_3_1_U19 ( .A1(Y1xD[13]), .A2(Y0xD[5]), .ZN(
        mul_y0y1_gf4_mul_3_1_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_3_1_U18 ( .A(mul_y0y1_gf4_mul_3_1_n75), .B(
        mul_y0y1_gf4_mul_3_1_n66), .Z(mul_y0y1_gf4_mul_3_1_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_1_U17 ( .A(mul_y0y1_gf4_mul_3_1_n65), .B(
        mul_y0y1_gf4_mul_3_1_n64), .ZN(mul_y0y1_gf4_mul_3_1_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_3_1_U16 ( .A1(mul_y0y1_gf4_mul_3_1_n63), .A2(
        mul_y0y1_gf4_mul_3_1_n62), .ZN(mul_y0y1_gf4_mul_3_1_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_1_U15 ( .A(mul_y0y1_gf4_mul_3_1_n61), .B(
        mul_y0y1_gf4_mul_3_1_n60), .ZN(mul_y0y1_gf4_mul_3_1_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_1_U14 ( .A(mul_y0y1_gf4_mul_3_1_n59), .B(
        mul_y0y1_gf4_mul_3_1_n58), .ZN(mul_y0y1_gf4_mul_3_1_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_1_U13 ( .A(mul_y0y1_gf4_mul_3_1_n57), .B(
        mul_y0y1_gf4_mul_3_1_n56), .ZN(mul_y0y1_Xi_mul_Yj_13__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_3_1_U12 ( .A1(Y1xD[12]), .A2(Y0xD[4]), .ZN(
        mul_y0y1_gf4_mul_3_1_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_3_1_U11 ( .A(mul_y0y1_gf4_mul_3_1_n66), .B(
        mul_y0y1_gf4_mul_3_1_n71), .Z(mul_y0y1_gf4_mul_3_1_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_1_U10 ( .A(mul_y0y1_gf4_mul_3_1_n55), .B(
        mul_y0y1_gf4_mul_3_1_n65), .ZN(mul_y0y1_gf4_mul_3_1_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_3_1_U9 ( .A1(mul_y0y1_gf4_mul_3_1_n61), .A2(
        mul_y0y1_gf4_mul_3_1_n59), .ZN(mul_y0y1_gf4_mul_3_1_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_1_U8 ( .A(Y1xD[12]), .B(Y1xD[14]), .ZN(
        mul_y0y1_gf4_mul_3_1_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_1_U7 ( .A(Y0xD[4]), .B(Y0xD[6]), .ZN(
        mul_y0y1_gf4_mul_3_1_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_3_1_U6 ( .A1(mul_y0y1_gf4_mul_3_1_n58), .A2(
        mul_y0y1_gf4_mul_3_1_n60), .ZN(mul_y0y1_gf4_mul_3_1_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_3_1_U5 ( .A(Y0xD[5]), .B(Y0xD[7]), .Z(
        mul_y0y1_gf4_mul_3_1_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_3_1_U4 ( .A(Y1xD[13]), .B(Y1xD[15]), .Z(
        mul_y0y1_gf4_mul_3_1_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_3_1_U3 ( .A1(mul_y0y1_gf4_mul_3_1_n54), .A2(
        mul_y0y1_gf4_mul_3_1_n53), .ZN(mul_y0y1_gf4_mul_3_1_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_1_U2 ( .A(Y1xD[12]), .B(Y1xD[13]), .ZN(
        mul_y0y1_gf4_mul_3_1_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_1_U1 ( .A(Y0xD[4]), .B(Y0xD[5]), .ZN(
        mul_y0y1_gf4_mul_3_1_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_0_U29 ( .A(mul_y0y1_gf4_mul_3_0_n77), .B(
        mul_y0y1_gf4_mul_3_0_n76), .ZN(mul_y0y1_Xi_mul_Yj_12__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_3_0_U28 ( .A1(Y1xD[15]), .A2(Y0xD[3]), .ZN(
        mul_y0y1_gf4_mul_3_0_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_3_0_U27 ( .A(mul_y0y1_gf4_mul_3_0_n75), .B(
        mul_y0y1_gf4_mul_3_0_n74), .Z(mul_y0y1_gf4_mul_3_0_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_0_U26 ( .A(mul_y0y1_gf4_mul_3_0_n73), .B(
        mul_y0y1_gf4_mul_3_0_n72), .ZN(mul_y0y1_Xi_mul_Yj_12__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_3_0_U25 ( .A1(Y1xD[14]), .A2(Y0xD[2]), .ZN(
        mul_y0y1_gf4_mul_3_0_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_3_0_U24 ( .A(mul_y0y1_gf4_mul_3_0_n74), .B(
        mul_y0y1_gf4_mul_3_0_n71), .Z(mul_y0y1_gf4_mul_3_0_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_3_0_U23 ( .A1(mul_y0y1_gf4_mul_3_0_n70), .A2(
        mul_y0y1_gf4_mul_3_0_n69), .ZN(mul_y0y1_gf4_mul_3_0_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_0_U22 ( .A(Y1xD[14]), .B(Y1xD[15]), .ZN(
        mul_y0y1_gf4_mul_3_0_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_0_U21 ( .A(Y0xD[2]), .B(Y0xD[3]), .ZN(
        mul_y0y1_gf4_mul_3_0_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_0_U20 ( .A(mul_y0y1_gf4_mul_3_0_n68), .B(
        mul_y0y1_gf4_mul_3_0_n67), .ZN(mul_y0y1_Xi_mul_Yj_12__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_3_0_U19 ( .A1(Y1xD[13]), .A2(Y0xD[1]), .ZN(
        mul_y0y1_gf4_mul_3_0_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_3_0_U18 ( .A(mul_y0y1_gf4_mul_3_0_n75), .B(
        mul_y0y1_gf4_mul_3_0_n66), .Z(mul_y0y1_gf4_mul_3_0_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_0_U17 ( .A(mul_y0y1_gf4_mul_3_0_n65), .B(
        mul_y0y1_gf4_mul_3_0_n64), .ZN(mul_y0y1_gf4_mul_3_0_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_3_0_U16 ( .A1(mul_y0y1_gf4_mul_3_0_n63), .A2(
        mul_y0y1_gf4_mul_3_0_n62), .ZN(mul_y0y1_gf4_mul_3_0_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_0_U15 ( .A(mul_y0y1_gf4_mul_3_0_n61), .B(
        mul_y0y1_gf4_mul_3_0_n60), .ZN(mul_y0y1_gf4_mul_3_0_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_0_U14 ( .A(mul_y0y1_gf4_mul_3_0_n59), .B(
        mul_y0y1_gf4_mul_3_0_n58), .ZN(mul_y0y1_gf4_mul_3_0_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_0_U13 ( .A(mul_y0y1_gf4_mul_3_0_n57), .B(
        mul_y0y1_gf4_mul_3_0_n56), .ZN(mul_y0y1_Xi_mul_Yj_12__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_3_0_U12 ( .A1(Y1xD[12]), .A2(Y0xD[0]), .ZN(
        mul_y0y1_gf4_mul_3_0_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_3_0_U11 ( .A(mul_y0y1_gf4_mul_3_0_n66), .B(
        mul_y0y1_gf4_mul_3_0_n71), .Z(mul_y0y1_gf4_mul_3_0_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_0_U10 ( .A(mul_y0y1_gf4_mul_3_0_n55), .B(
        mul_y0y1_gf4_mul_3_0_n65), .ZN(mul_y0y1_gf4_mul_3_0_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_3_0_U9 ( .A1(mul_y0y1_gf4_mul_3_0_n61), .A2(
        mul_y0y1_gf4_mul_3_0_n59), .ZN(mul_y0y1_gf4_mul_3_0_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_0_U8 ( .A(Y1xD[12]), .B(Y1xD[14]), .ZN(
        mul_y0y1_gf4_mul_3_0_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_0_U7 ( .A(Y0xD[0]), .B(Y0xD[2]), .ZN(
        mul_y0y1_gf4_mul_3_0_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_3_0_U6 ( .A1(mul_y0y1_gf4_mul_3_0_n58), .A2(
        mul_y0y1_gf4_mul_3_0_n60), .ZN(mul_y0y1_gf4_mul_3_0_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_3_0_U5 ( .A(Y0xD[1]), .B(Y0xD[3]), .Z(
        mul_y0y1_gf4_mul_3_0_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_3_0_U4 ( .A(Y1xD[13]), .B(Y1xD[15]), .Z(
        mul_y0y1_gf4_mul_3_0_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_3_0_U3 ( .A1(mul_y0y1_gf4_mul_3_0_n54), .A2(
        mul_y0y1_gf4_mul_3_0_n53), .ZN(mul_y0y1_gf4_mul_3_0_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_0_U2 ( .A(Y1xD[12]), .B(Y1xD[13]), .ZN(
        mul_y0y1_gf4_mul_3_0_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_3_0_U1 ( .A(Y0xD[0]), .B(Y0xD[1]), .ZN(
        mul_y0y1_gf4_mul_3_0_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_3_U29 ( .A(mul_y0y1_gf4_mul_2_3_n77), .B(
        mul_y0y1_gf4_mul_2_3_n76), .ZN(mul_y0y1_Xi_mul_Yj_11__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_3_U28 ( .A1(Y1xD[11]), .A2(Y0xD[15]), .ZN(
        mul_y0y1_gf4_mul_2_3_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_2_3_U27 ( .A(mul_y0y1_gf4_mul_2_3_n75), .B(
        mul_y0y1_gf4_mul_2_3_n74), .Z(mul_y0y1_gf4_mul_2_3_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_3_U26 ( .A(mul_y0y1_gf4_mul_2_3_n73), .B(
        mul_y0y1_gf4_mul_2_3_n72), .ZN(mul_y0y1_Xi_mul_Yj_11__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_3_U25 ( .A1(Y1xD[10]), .A2(Y0xD[14]), .ZN(
        mul_y0y1_gf4_mul_2_3_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_2_3_U24 ( .A(mul_y0y1_gf4_mul_2_3_n74), .B(
        mul_y0y1_gf4_mul_2_3_n71), .Z(mul_y0y1_gf4_mul_2_3_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_2_3_U23 ( .A1(mul_y0y1_gf4_mul_2_3_n70), .A2(
        mul_y0y1_gf4_mul_2_3_n69), .ZN(mul_y0y1_gf4_mul_2_3_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_3_U22 ( .A(Y1xD[10]), .B(Y1xD[11]), .ZN(
        mul_y0y1_gf4_mul_2_3_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_3_U21 ( .A(Y0xD[14]), .B(Y0xD[15]), .ZN(
        mul_y0y1_gf4_mul_2_3_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_3_U20 ( .A(mul_y0y1_gf4_mul_2_3_n68), .B(
        mul_y0y1_gf4_mul_2_3_n67), .ZN(mul_y0y1_Xi_mul_Yj_11__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_3_U19 ( .A1(Y1xD[9]), .A2(Y0xD[13]), .ZN(
        mul_y0y1_gf4_mul_2_3_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_2_3_U18 ( .A(mul_y0y1_gf4_mul_2_3_n75), .B(
        mul_y0y1_gf4_mul_2_3_n66), .Z(mul_y0y1_gf4_mul_2_3_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_3_U17 ( .A(mul_y0y1_gf4_mul_2_3_n65), .B(
        mul_y0y1_gf4_mul_2_3_n64), .ZN(mul_y0y1_gf4_mul_2_3_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_2_3_U16 ( .A1(mul_y0y1_gf4_mul_2_3_n63), .A2(
        mul_y0y1_gf4_mul_2_3_n62), .ZN(mul_y0y1_gf4_mul_2_3_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_3_U15 ( .A(mul_y0y1_gf4_mul_2_3_n61), .B(
        mul_y0y1_gf4_mul_2_3_n60), .ZN(mul_y0y1_gf4_mul_2_3_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_3_U14 ( .A(mul_y0y1_gf4_mul_2_3_n59), .B(
        mul_y0y1_gf4_mul_2_3_n58), .ZN(mul_y0y1_gf4_mul_2_3_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_3_U13 ( .A(mul_y0y1_gf4_mul_2_3_n57), .B(
        mul_y0y1_gf4_mul_2_3_n56), .ZN(mul_y0y1_Xi_mul_Yj_11__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_3_U12 ( .A1(Y1xD[8]), .A2(Y0xD[12]), .ZN(
        mul_y0y1_gf4_mul_2_3_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_2_3_U11 ( .A(mul_y0y1_gf4_mul_2_3_n66), .B(
        mul_y0y1_gf4_mul_2_3_n71), .Z(mul_y0y1_gf4_mul_2_3_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_3_U10 ( .A(mul_y0y1_gf4_mul_2_3_n55), .B(
        mul_y0y1_gf4_mul_2_3_n65), .ZN(mul_y0y1_gf4_mul_2_3_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_2_3_U9 ( .A1(mul_y0y1_gf4_mul_2_3_n61), .A2(
        mul_y0y1_gf4_mul_2_3_n59), .ZN(mul_y0y1_gf4_mul_2_3_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_3_U8 ( .A(Y1xD[8]), .B(Y1xD[10]), .ZN(
        mul_y0y1_gf4_mul_2_3_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_3_U7 ( .A(Y0xD[12]), .B(Y0xD[14]), .ZN(
        mul_y0y1_gf4_mul_2_3_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_2_3_U6 ( .A1(mul_y0y1_gf4_mul_2_3_n58), .A2(
        mul_y0y1_gf4_mul_2_3_n60), .ZN(mul_y0y1_gf4_mul_2_3_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_2_3_U5 ( .A(Y0xD[13]), .B(Y0xD[15]), .Z(
        mul_y0y1_gf4_mul_2_3_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_2_3_U4 ( .A(Y1xD[9]), .B(Y1xD[11]), .Z(
        mul_y0y1_gf4_mul_2_3_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_2_3_U3 ( .A1(mul_y0y1_gf4_mul_2_3_n54), .A2(
        mul_y0y1_gf4_mul_2_3_n53), .ZN(mul_y0y1_gf4_mul_2_3_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_3_U2 ( .A(Y1xD[8]), .B(Y1xD[9]), .ZN(
        mul_y0y1_gf4_mul_2_3_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_3_U1 ( .A(Y0xD[12]), .B(Y0xD[13]), .ZN(
        mul_y0y1_gf4_mul_2_3_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U29 ( .A(mul_y0y1_gf4_mul_2_2_n77), .B(
        mul_y0y1_gf4_mul_2_2_n76), .ZN(mul_y0y1_FFxDN[43]) );
  NAND2_X1 mul_y0y1_gf4_mul_2_2_U28 ( .A1(Y1xD[11]), .A2(Y0xD[11]), .ZN(
        mul_y0y1_gf4_mul_2_2_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_2_2_U27 ( .A(mul_y0y1_gf4_mul_2_2_n75), .B(
        mul_y0y1_gf4_mul_2_2_n74), .Z(mul_y0y1_gf4_mul_2_2_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U26 ( .A(mul_y0y1_gf4_mul_2_2_n73), .B(
        mul_y0y1_gf4_mul_2_2_n72), .ZN(mul_y0y1_FFxDN[42]) );
  NAND2_X1 mul_y0y1_gf4_mul_2_2_U25 ( .A1(Y1xD[10]), .A2(Y0xD[10]), .ZN(
        mul_y0y1_gf4_mul_2_2_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_2_2_U24 ( .A(mul_y0y1_gf4_mul_2_2_n74), .B(
        mul_y0y1_gf4_mul_2_2_n71), .Z(mul_y0y1_gf4_mul_2_2_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_2_2_U23 ( .A1(mul_y0y1_gf4_mul_2_2_n70), .A2(
        mul_y0y1_gf4_mul_2_2_n69), .ZN(mul_y0y1_gf4_mul_2_2_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U22 ( .A(Y1xD[10]), .B(Y1xD[11]), .ZN(
        mul_y0y1_gf4_mul_2_2_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U21 ( .A(Y0xD[10]), .B(Y0xD[11]), .ZN(
        mul_y0y1_gf4_mul_2_2_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U20 ( .A(mul_y0y1_gf4_mul_2_2_n68), .B(
        mul_y0y1_gf4_mul_2_2_n67), .ZN(mul_y0y1_FFxDN[41]) );
  NAND2_X1 mul_y0y1_gf4_mul_2_2_U19 ( .A1(Y1xD[9]), .A2(Y0xD[9]), .ZN(
        mul_y0y1_gf4_mul_2_2_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_2_2_U18 ( .A(mul_y0y1_gf4_mul_2_2_n75), .B(
        mul_y0y1_gf4_mul_2_2_n66), .Z(mul_y0y1_gf4_mul_2_2_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U17 ( .A(mul_y0y1_gf4_mul_2_2_n65), .B(
        mul_y0y1_gf4_mul_2_2_n64), .ZN(mul_y0y1_gf4_mul_2_2_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_2_2_U16 ( .A1(mul_y0y1_gf4_mul_2_2_n63), .A2(
        mul_y0y1_gf4_mul_2_2_n62), .ZN(mul_y0y1_gf4_mul_2_2_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U15 ( .A(mul_y0y1_gf4_mul_2_2_n61), .B(
        mul_y0y1_gf4_mul_2_2_n60), .ZN(mul_y0y1_gf4_mul_2_2_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U14 ( .A(mul_y0y1_gf4_mul_2_2_n59), .B(
        mul_y0y1_gf4_mul_2_2_n58), .ZN(mul_y0y1_gf4_mul_2_2_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U13 ( .A(mul_y0y1_gf4_mul_2_2_n57), .B(
        mul_y0y1_gf4_mul_2_2_n56), .ZN(mul_y0y1_FFxDN[40]) );
  NAND2_X1 mul_y0y1_gf4_mul_2_2_U12 ( .A1(Y1xD[8]), .A2(Y0xD[8]), .ZN(
        mul_y0y1_gf4_mul_2_2_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_2_2_U11 ( .A(mul_y0y1_gf4_mul_2_2_n66), .B(
        mul_y0y1_gf4_mul_2_2_n71), .Z(mul_y0y1_gf4_mul_2_2_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U10 ( .A(mul_y0y1_gf4_mul_2_2_n55), .B(
        mul_y0y1_gf4_mul_2_2_n65), .ZN(mul_y0y1_gf4_mul_2_2_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_2_2_U9 ( .A1(mul_y0y1_gf4_mul_2_2_n61), .A2(
        mul_y0y1_gf4_mul_2_2_n59), .ZN(mul_y0y1_gf4_mul_2_2_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U8 ( .A(Y1xD[8]), .B(Y1xD[10]), .ZN(
        mul_y0y1_gf4_mul_2_2_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U7 ( .A(Y0xD[8]), .B(Y0xD[10]), .ZN(
        mul_y0y1_gf4_mul_2_2_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_2_2_U6 ( .A1(mul_y0y1_gf4_mul_2_2_n58), .A2(
        mul_y0y1_gf4_mul_2_2_n60), .ZN(mul_y0y1_gf4_mul_2_2_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_2_2_U5 ( .A(Y0xD[9]), .B(Y0xD[11]), .Z(
        mul_y0y1_gf4_mul_2_2_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_2_2_U4 ( .A(Y1xD[9]), .B(Y1xD[11]), .Z(
        mul_y0y1_gf4_mul_2_2_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_2_2_U3 ( .A1(mul_y0y1_gf4_mul_2_2_n54), .A2(
        mul_y0y1_gf4_mul_2_2_n53), .ZN(mul_y0y1_gf4_mul_2_2_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U2 ( .A(Y1xD[8]), .B(Y1xD[9]), .ZN(
        mul_y0y1_gf4_mul_2_2_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_2_U1 ( .A(Y0xD[8]), .B(Y0xD[9]), .ZN(
        mul_y0y1_gf4_mul_2_2_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U29 ( .A(mul_y0y1_gf4_mul_2_1_n77), .B(
        mul_y0y1_gf4_mul_2_1_n76), .ZN(mul_y0y1_Xi_mul_Yj_9__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_1_U28 ( .A1(Y1xD[11]), .A2(Y0xD[7]), .ZN(
        mul_y0y1_gf4_mul_2_1_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_2_1_U27 ( .A(mul_y0y1_gf4_mul_2_1_n75), .B(
        mul_y0y1_gf4_mul_2_1_n74), .Z(mul_y0y1_gf4_mul_2_1_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U26 ( .A(mul_y0y1_gf4_mul_2_1_n73), .B(
        mul_y0y1_gf4_mul_2_1_n72), .ZN(mul_y0y1_Xi_mul_Yj_9__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_1_U25 ( .A1(Y1xD[10]), .A2(Y0xD[6]), .ZN(
        mul_y0y1_gf4_mul_2_1_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_2_1_U24 ( .A(mul_y0y1_gf4_mul_2_1_n74), .B(
        mul_y0y1_gf4_mul_2_1_n71), .Z(mul_y0y1_gf4_mul_2_1_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_2_1_U23 ( .A1(mul_y0y1_gf4_mul_2_1_n70), .A2(
        mul_y0y1_gf4_mul_2_1_n69), .ZN(mul_y0y1_gf4_mul_2_1_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U22 ( .A(Y1xD[10]), .B(Y1xD[11]), .ZN(
        mul_y0y1_gf4_mul_2_1_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U21 ( .A(Y0xD[6]), .B(Y0xD[7]), .ZN(
        mul_y0y1_gf4_mul_2_1_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U20 ( .A(mul_y0y1_gf4_mul_2_1_n68), .B(
        mul_y0y1_gf4_mul_2_1_n67), .ZN(mul_y0y1_Xi_mul_Yj_9__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_1_U19 ( .A1(Y1xD[9]), .A2(Y0xD[5]), .ZN(
        mul_y0y1_gf4_mul_2_1_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_2_1_U18 ( .A(mul_y0y1_gf4_mul_2_1_n75), .B(
        mul_y0y1_gf4_mul_2_1_n66), .Z(mul_y0y1_gf4_mul_2_1_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U17 ( .A(mul_y0y1_gf4_mul_2_1_n65), .B(
        mul_y0y1_gf4_mul_2_1_n64), .ZN(mul_y0y1_gf4_mul_2_1_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_2_1_U16 ( .A1(mul_y0y1_gf4_mul_2_1_n63), .A2(
        mul_y0y1_gf4_mul_2_1_n62), .ZN(mul_y0y1_gf4_mul_2_1_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U15 ( .A(mul_y0y1_gf4_mul_2_1_n61), .B(
        mul_y0y1_gf4_mul_2_1_n60), .ZN(mul_y0y1_gf4_mul_2_1_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U14 ( .A(mul_y0y1_gf4_mul_2_1_n59), .B(
        mul_y0y1_gf4_mul_2_1_n58), .ZN(mul_y0y1_gf4_mul_2_1_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U13 ( .A(mul_y0y1_gf4_mul_2_1_n57), .B(
        mul_y0y1_gf4_mul_2_1_n56), .ZN(mul_y0y1_Xi_mul_Yj_9__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_1_U12 ( .A1(Y1xD[8]), .A2(Y0xD[4]), .ZN(
        mul_y0y1_gf4_mul_2_1_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_2_1_U11 ( .A(mul_y0y1_gf4_mul_2_1_n66), .B(
        mul_y0y1_gf4_mul_2_1_n71), .Z(mul_y0y1_gf4_mul_2_1_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U10 ( .A(mul_y0y1_gf4_mul_2_1_n55), .B(
        mul_y0y1_gf4_mul_2_1_n65), .ZN(mul_y0y1_gf4_mul_2_1_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_2_1_U9 ( .A1(mul_y0y1_gf4_mul_2_1_n61), .A2(
        mul_y0y1_gf4_mul_2_1_n59), .ZN(mul_y0y1_gf4_mul_2_1_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U8 ( .A(Y1xD[8]), .B(Y1xD[10]), .ZN(
        mul_y0y1_gf4_mul_2_1_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U7 ( .A(Y0xD[4]), .B(Y0xD[6]), .ZN(
        mul_y0y1_gf4_mul_2_1_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_2_1_U6 ( .A1(mul_y0y1_gf4_mul_2_1_n58), .A2(
        mul_y0y1_gf4_mul_2_1_n60), .ZN(mul_y0y1_gf4_mul_2_1_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_2_1_U5 ( .A(Y0xD[5]), .B(Y0xD[7]), .Z(
        mul_y0y1_gf4_mul_2_1_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_2_1_U4 ( .A(Y1xD[9]), .B(Y1xD[11]), .Z(
        mul_y0y1_gf4_mul_2_1_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_2_1_U3 ( .A1(mul_y0y1_gf4_mul_2_1_n54), .A2(
        mul_y0y1_gf4_mul_2_1_n53), .ZN(mul_y0y1_gf4_mul_2_1_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U2 ( .A(Y1xD[8]), .B(Y1xD[9]), .ZN(
        mul_y0y1_gf4_mul_2_1_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_1_U1 ( .A(Y0xD[4]), .B(Y0xD[5]), .ZN(
        mul_y0y1_gf4_mul_2_1_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U29 ( .A(mul_y0y1_gf4_mul_2_0_n77), .B(
        mul_y0y1_gf4_mul_2_0_n76), .ZN(mul_y0y1_Xi_mul_Yj_8__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_0_U28 ( .A1(Y1xD[11]), .A2(Y0xD[3]), .ZN(
        mul_y0y1_gf4_mul_2_0_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_2_0_U27 ( .A(mul_y0y1_gf4_mul_2_0_n75), .B(
        mul_y0y1_gf4_mul_2_0_n74), .Z(mul_y0y1_gf4_mul_2_0_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U26 ( .A(mul_y0y1_gf4_mul_2_0_n73), .B(
        mul_y0y1_gf4_mul_2_0_n72), .ZN(mul_y0y1_Xi_mul_Yj_8__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_0_U25 ( .A1(Y1xD[10]), .A2(Y0xD[2]), .ZN(
        mul_y0y1_gf4_mul_2_0_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_2_0_U24 ( .A(mul_y0y1_gf4_mul_2_0_n74), .B(
        mul_y0y1_gf4_mul_2_0_n71), .Z(mul_y0y1_gf4_mul_2_0_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_2_0_U23 ( .A1(mul_y0y1_gf4_mul_2_0_n70), .A2(
        mul_y0y1_gf4_mul_2_0_n69), .ZN(mul_y0y1_gf4_mul_2_0_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U22 ( .A(Y1xD[10]), .B(Y1xD[11]), .ZN(
        mul_y0y1_gf4_mul_2_0_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U21 ( .A(Y0xD[2]), .B(Y0xD[3]), .ZN(
        mul_y0y1_gf4_mul_2_0_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U20 ( .A(mul_y0y1_gf4_mul_2_0_n68), .B(
        mul_y0y1_gf4_mul_2_0_n67), .ZN(mul_y0y1_Xi_mul_Yj_8__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_0_U19 ( .A1(Y1xD[9]), .A2(Y0xD[1]), .ZN(
        mul_y0y1_gf4_mul_2_0_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_2_0_U18 ( .A(mul_y0y1_gf4_mul_2_0_n75), .B(
        mul_y0y1_gf4_mul_2_0_n66), .Z(mul_y0y1_gf4_mul_2_0_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U17 ( .A(mul_y0y1_gf4_mul_2_0_n65), .B(
        mul_y0y1_gf4_mul_2_0_n64), .ZN(mul_y0y1_gf4_mul_2_0_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_2_0_U16 ( .A1(mul_y0y1_gf4_mul_2_0_n63), .A2(
        mul_y0y1_gf4_mul_2_0_n62), .ZN(mul_y0y1_gf4_mul_2_0_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U15 ( .A(mul_y0y1_gf4_mul_2_0_n61), .B(
        mul_y0y1_gf4_mul_2_0_n60), .ZN(mul_y0y1_gf4_mul_2_0_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U14 ( .A(mul_y0y1_gf4_mul_2_0_n59), .B(
        mul_y0y1_gf4_mul_2_0_n58), .ZN(mul_y0y1_gf4_mul_2_0_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U13 ( .A(mul_y0y1_gf4_mul_2_0_n57), .B(
        mul_y0y1_gf4_mul_2_0_n56), .ZN(mul_y0y1_Xi_mul_Yj_8__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_2_0_U12 ( .A1(Y1xD[8]), .A2(Y0xD[0]), .ZN(
        mul_y0y1_gf4_mul_2_0_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_2_0_U11 ( .A(mul_y0y1_gf4_mul_2_0_n66), .B(
        mul_y0y1_gf4_mul_2_0_n71), .Z(mul_y0y1_gf4_mul_2_0_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U10 ( .A(mul_y0y1_gf4_mul_2_0_n55), .B(
        mul_y0y1_gf4_mul_2_0_n65), .ZN(mul_y0y1_gf4_mul_2_0_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_2_0_U9 ( .A1(mul_y0y1_gf4_mul_2_0_n61), .A2(
        mul_y0y1_gf4_mul_2_0_n59), .ZN(mul_y0y1_gf4_mul_2_0_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U8 ( .A(Y1xD[8]), .B(Y1xD[10]), .ZN(
        mul_y0y1_gf4_mul_2_0_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U7 ( .A(Y0xD[0]), .B(Y0xD[2]), .ZN(
        mul_y0y1_gf4_mul_2_0_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_2_0_U6 ( .A1(mul_y0y1_gf4_mul_2_0_n58), .A2(
        mul_y0y1_gf4_mul_2_0_n60), .ZN(mul_y0y1_gf4_mul_2_0_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_2_0_U5 ( .A(Y0xD[1]), .B(Y0xD[3]), .Z(
        mul_y0y1_gf4_mul_2_0_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_2_0_U4 ( .A(Y1xD[9]), .B(Y1xD[11]), .Z(
        mul_y0y1_gf4_mul_2_0_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_2_0_U3 ( .A1(mul_y0y1_gf4_mul_2_0_n54), .A2(
        mul_y0y1_gf4_mul_2_0_n53), .ZN(mul_y0y1_gf4_mul_2_0_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U2 ( .A(Y1xD[8]), .B(Y1xD[9]), .ZN(
        mul_y0y1_gf4_mul_2_0_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_2_0_U1 ( .A(Y0xD[0]), .B(Y0xD[1]), .ZN(
        mul_y0y1_gf4_mul_2_0_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_3_U29 ( .A(mul_y0y1_gf4_mul_1_3_n77), .B(
        mul_y0y1_gf4_mul_1_3_n76), .ZN(mul_y0y1_Xi_mul_Yj_7__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_3_U28 ( .A1(Y1xD[7]), .A2(Y0xD[15]), .ZN(
        mul_y0y1_gf4_mul_1_3_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_1_3_U27 ( .A(mul_y0y1_gf4_mul_1_3_n75), .B(
        mul_y0y1_gf4_mul_1_3_n74), .Z(mul_y0y1_gf4_mul_1_3_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_3_U26 ( .A(mul_y0y1_gf4_mul_1_3_n73), .B(
        mul_y0y1_gf4_mul_1_3_n72), .ZN(mul_y0y1_Xi_mul_Yj_7__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_3_U25 ( .A1(Y1xD[6]), .A2(Y0xD[14]), .ZN(
        mul_y0y1_gf4_mul_1_3_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_1_3_U24 ( .A(mul_y0y1_gf4_mul_1_3_n74), .B(
        mul_y0y1_gf4_mul_1_3_n71), .Z(mul_y0y1_gf4_mul_1_3_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_1_3_U23 ( .A1(mul_y0y1_gf4_mul_1_3_n70), .A2(
        mul_y0y1_gf4_mul_1_3_n69), .ZN(mul_y0y1_gf4_mul_1_3_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_3_U22 ( .A(Y1xD[6]), .B(Y1xD[7]), .ZN(
        mul_y0y1_gf4_mul_1_3_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_3_U21 ( .A(Y0xD[14]), .B(Y0xD[15]), .ZN(
        mul_y0y1_gf4_mul_1_3_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_3_U20 ( .A(mul_y0y1_gf4_mul_1_3_n68), .B(
        mul_y0y1_gf4_mul_1_3_n67), .ZN(mul_y0y1_Xi_mul_Yj_7__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_3_U19 ( .A1(Y1xD[5]), .A2(Y0xD[13]), .ZN(
        mul_y0y1_gf4_mul_1_3_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_1_3_U18 ( .A(mul_y0y1_gf4_mul_1_3_n75), .B(
        mul_y0y1_gf4_mul_1_3_n66), .Z(mul_y0y1_gf4_mul_1_3_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_3_U17 ( .A(mul_y0y1_gf4_mul_1_3_n65), .B(
        mul_y0y1_gf4_mul_1_3_n64), .ZN(mul_y0y1_gf4_mul_1_3_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_1_3_U16 ( .A1(mul_y0y1_gf4_mul_1_3_n63), .A2(
        mul_y0y1_gf4_mul_1_3_n62), .ZN(mul_y0y1_gf4_mul_1_3_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_3_U15 ( .A(mul_y0y1_gf4_mul_1_3_n61), .B(
        mul_y0y1_gf4_mul_1_3_n60), .ZN(mul_y0y1_gf4_mul_1_3_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_3_U14 ( .A(mul_y0y1_gf4_mul_1_3_n59), .B(
        mul_y0y1_gf4_mul_1_3_n58), .ZN(mul_y0y1_gf4_mul_1_3_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_3_U13 ( .A(mul_y0y1_gf4_mul_1_3_n57), .B(
        mul_y0y1_gf4_mul_1_3_n56), .ZN(mul_y0y1_Xi_mul_Yj_7__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_3_U12 ( .A1(Y1xD[4]), .A2(Y0xD[12]), .ZN(
        mul_y0y1_gf4_mul_1_3_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_1_3_U11 ( .A(mul_y0y1_gf4_mul_1_3_n66), .B(
        mul_y0y1_gf4_mul_1_3_n71), .Z(mul_y0y1_gf4_mul_1_3_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_3_U10 ( .A(mul_y0y1_gf4_mul_1_3_n55), .B(
        mul_y0y1_gf4_mul_1_3_n65), .ZN(mul_y0y1_gf4_mul_1_3_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_1_3_U9 ( .A1(mul_y0y1_gf4_mul_1_3_n61), .A2(
        mul_y0y1_gf4_mul_1_3_n59), .ZN(mul_y0y1_gf4_mul_1_3_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_3_U8 ( .A(Y1xD[4]), .B(Y1xD[6]), .ZN(
        mul_y0y1_gf4_mul_1_3_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_3_U7 ( .A(Y0xD[12]), .B(Y0xD[14]), .ZN(
        mul_y0y1_gf4_mul_1_3_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_1_3_U6 ( .A1(mul_y0y1_gf4_mul_1_3_n58), .A2(
        mul_y0y1_gf4_mul_1_3_n60), .ZN(mul_y0y1_gf4_mul_1_3_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_1_3_U5 ( .A(Y0xD[13]), .B(Y0xD[15]), .Z(
        mul_y0y1_gf4_mul_1_3_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_1_3_U4 ( .A(Y1xD[5]), .B(Y1xD[7]), .Z(
        mul_y0y1_gf4_mul_1_3_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_1_3_U3 ( .A1(mul_y0y1_gf4_mul_1_3_n54), .A2(
        mul_y0y1_gf4_mul_1_3_n53), .ZN(mul_y0y1_gf4_mul_1_3_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_3_U2 ( .A(Y1xD[4]), .B(Y1xD[5]), .ZN(
        mul_y0y1_gf4_mul_1_3_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_3_U1 ( .A(Y0xD[12]), .B(Y0xD[13]), .ZN(
        mul_y0y1_gf4_mul_1_3_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U29 ( .A(mul_y0y1_gf4_mul_1_2_n77), .B(
        mul_y0y1_gf4_mul_1_2_n76), .ZN(mul_y0y1_Xi_mul_Yj_6__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_2_U28 ( .A1(Y1xD[7]), .A2(Y0xD[11]), .ZN(
        mul_y0y1_gf4_mul_1_2_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_1_2_U27 ( .A(mul_y0y1_gf4_mul_1_2_n75), .B(
        mul_y0y1_gf4_mul_1_2_n74), .Z(mul_y0y1_gf4_mul_1_2_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U26 ( .A(mul_y0y1_gf4_mul_1_2_n73), .B(
        mul_y0y1_gf4_mul_1_2_n72), .ZN(mul_y0y1_Xi_mul_Yj_6__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_2_U25 ( .A1(Y1xD[6]), .A2(Y0xD[10]), .ZN(
        mul_y0y1_gf4_mul_1_2_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_1_2_U24 ( .A(mul_y0y1_gf4_mul_1_2_n74), .B(
        mul_y0y1_gf4_mul_1_2_n71), .Z(mul_y0y1_gf4_mul_1_2_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_1_2_U23 ( .A1(mul_y0y1_gf4_mul_1_2_n70), .A2(
        mul_y0y1_gf4_mul_1_2_n69), .ZN(mul_y0y1_gf4_mul_1_2_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U22 ( .A(Y1xD[6]), .B(Y1xD[7]), .ZN(
        mul_y0y1_gf4_mul_1_2_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U21 ( .A(Y0xD[10]), .B(Y0xD[11]), .ZN(
        mul_y0y1_gf4_mul_1_2_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U20 ( .A(mul_y0y1_gf4_mul_1_2_n68), .B(
        mul_y0y1_gf4_mul_1_2_n67), .ZN(mul_y0y1_Xi_mul_Yj_6__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_2_U19 ( .A1(Y1xD[5]), .A2(Y0xD[9]), .ZN(
        mul_y0y1_gf4_mul_1_2_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_1_2_U18 ( .A(mul_y0y1_gf4_mul_1_2_n75), .B(
        mul_y0y1_gf4_mul_1_2_n66), .Z(mul_y0y1_gf4_mul_1_2_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U17 ( .A(mul_y0y1_gf4_mul_1_2_n65), .B(
        mul_y0y1_gf4_mul_1_2_n64), .ZN(mul_y0y1_gf4_mul_1_2_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_1_2_U16 ( .A1(mul_y0y1_gf4_mul_1_2_n63), .A2(
        mul_y0y1_gf4_mul_1_2_n62), .ZN(mul_y0y1_gf4_mul_1_2_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U15 ( .A(mul_y0y1_gf4_mul_1_2_n61), .B(
        mul_y0y1_gf4_mul_1_2_n60), .ZN(mul_y0y1_gf4_mul_1_2_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U14 ( .A(mul_y0y1_gf4_mul_1_2_n59), .B(
        mul_y0y1_gf4_mul_1_2_n58), .ZN(mul_y0y1_gf4_mul_1_2_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U13 ( .A(mul_y0y1_gf4_mul_1_2_n57), .B(
        mul_y0y1_gf4_mul_1_2_n56), .ZN(mul_y0y1_Xi_mul_Yj_6__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_2_U12 ( .A1(Y1xD[4]), .A2(Y0xD[8]), .ZN(
        mul_y0y1_gf4_mul_1_2_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_1_2_U11 ( .A(mul_y0y1_gf4_mul_1_2_n66), .B(
        mul_y0y1_gf4_mul_1_2_n71), .Z(mul_y0y1_gf4_mul_1_2_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U10 ( .A(mul_y0y1_gf4_mul_1_2_n55), .B(
        mul_y0y1_gf4_mul_1_2_n65), .ZN(mul_y0y1_gf4_mul_1_2_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_1_2_U9 ( .A1(mul_y0y1_gf4_mul_1_2_n61), .A2(
        mul_y0y1_gf4_mul_1_2_n59), .ZN(mul_y0y1_gf4_mul_1_2_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U8 ( .A(Y1xD[4]), .B(Y1xD[6]), .ZN(
        mul_y0y1_gf4_mul_1_2_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U7 ( .A(Y0xD[8]), .B(Y0xD[10]), .ZN(
        mul_y0y1_gf4_mul_1_2_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_1_2_U6 ( .A1(mul_y0y1_gf4_mul_1_2_n58), .A2(
        mul_y0y1_gf4_mul_1_2_n60), .ZN(mul_y0y1_gf4_mul_1_2_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_1_2_U5 ( .A(Y0xD[9]), .B(Y0xD[11]), .Z(
        mul_y0y1_gf4_mul_1_2_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_1_2_U4 ( .A(Y1xD[5]), .B(Y1xD[7]), .Z(
        mul_y0y1_gf4_mul_1_2_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_1_2_U3 ( .A1(mul_y0y1_gf4_mul_1_2_n54), .A2(
        mul_y0y1_gf4_mul_1_2_n53), .ZN(mul_y0y1_gf4_mul_1_2_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U2 ( .A(Y1xD[4]), .B(Y1xD[5]), .ZN(
        mul_y0y1_gf4_mul_1_2_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_2_U1 ( .A(Y0xD[8]), .B(Y0xD[9]), .ZN(
        mul_y0y1_gf4_mul_1_2_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U29 ( .A(mul_y0y1_gf4_mul_1_1_n77), .B(
        mul_y0y1_gf4_mul_1_1_n76), .ZN(mul_y0y1_FFxDN[23]) );
  NAND2_X1 mul_y0y1_gf4_mul_1_1_U28 ( .A1(Y1xD[7]), .A2(Y0xD[7]), .ZN(
        mul_y0y1_gf4_mul_1_1_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_1_1_U27 ( .A(mul_y0y1_gf4_mul_1_1_n75), .B(
        mul_y0y1_gf4_mul_1_1_n74), .Z(mul_y0y1_gf4_mul_1_1_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U26 ( .A(mul_y0y1_gf4_mul_1_1_n73), .B(
        mul_y0y1_gf4_mul_1_1_n72), .ZN(mul_y0y1_FFxDN[22]) );
  NAND2_X1 mul_y0y1_gf4_mul_1_1_U25 ( .A1(Y1xD[6]), .A2(Y0xD[6]), .ZN(
        mul_y0y1_gf4_mul_1_1_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_1_1_U24 ( .A(mul_y0y1_gf4_mul_1_1_n74), .B(
        mul_y0y1_gf4_mul_1_1_n71), .Z(mul_y0y1_gf4_mul_1_1_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_1_1_U23 ( .A1(mul_y0y1_gf4_mul_1_1_n70), .A2(
        mul_y0y1_gf4_mul_1_1_n69), .ZN(mul_y0y1_gf4_mul_1_1_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U22 ( .A(Y1xD[6]), .B(Y1xD[7]), .ZN(
        mul_y0y1_gf4_mul_1_1_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U21 ( .A(Y0xD[6]), .B(Y0xD[7]), .ZN(
        mul_y0y1_gf4_mul_1_1_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U20 ( .A(mul_y0y1_gf4_mul_1_1_n68), .B(
        mul_y0y1_gf4_mul_1_1_n67), .ZN(mul_y0y1_FFxDN[21]) );
  NAND2_X1 mul_y0y1_gf4_mul_1_1_U19 ( .A1(Y1xD[5]), .A2(Y0xD[5]), .ZN(
        mul_y0y1_gf4_mul_1_1_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_1_1_U18 ( .A(mul_y0y1_gf4_mul_1_1_n75), .B(
        mul_y0y1_gf4_mul_1_1_n66), .Z(mul_y0y1_gf4_mul_1_1_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U17 ( .A(mul_y0y1_gf4_mul_1_1_n65), .B(
        mul_y0y1_gf4_mul_1_1_n64), .ZN(mul_y0y1_gf4_mul_1_1_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_1_1_U16 ( .A1(mul_y0y1_gf4_mul_1_1_n63), .A2(
        mul_y0y1_gf4_mul_1_1_n62), .ZN(mul_y0y1_gf4_mul_1_1_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U15 ( .A(mul_y0y1_gf4_mul_1_1_n61), .B(
        mul_y0y1_gf4_mul_1_1_n60), .ZN(mul_y0y1_gf4_mul_1_1_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U14 ( .A(mul_y0y1_gf4_mul_1_1_n59), .B(
        mul_y0y1_gf4_mul_1_1_n58), .ZN(mul_y0y1_gf4_mul_1_1_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U13 ( .A(mul_y0y1_gf4_mul_1_1_n57), .B(
        mul_y0y1_gf4_mul_1_1_n56), .ZN(mul_y0y1_FFxDN[20]) );
  NAND2_X1 mul_y0y1_gf4_mul_1_1_U12 ( .A1(Y1xD[4]), .A2(Y0xD[4]), .ZN(
        mul_y0y1_gf4_mul_1_1_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_1_1_U11 ( .A(mul_y0y1_gf4_mul_1_1_n66), .B(
        mul_y0y1_gf4_mul_1_1_n71), .Z(mul_y0y1_gf4_mul_1_1_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U10 ( .A(mul_y0y1_gf4_mul_1_1_n55), .B(
        mul_y0y1_gf4_mul_1_1_n65), .ZN(mul_y0y1_gf4_mul_1_1_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_1_1_U9 ( .A1(mul_y0y1_gf4_mul_1_1_n61), .A2(
        mul_y0y1_gf4_mul_1_1_n59), .ZN(mul_y0y1_gf4_mul_1_1_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U8 ( .A(Y1xD[4]), .B(Y1xD[6]), .ZN(
        mul_y0y1_gf4_mul_1_1_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U7 ( .A(Y0xD[4]), .B(Y0xD[6]), .ZN(
        mul_y0y1_gf4_mul_1_1_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_1_1_U6 ( .A1(mul_y0y1_gf4_mul_1_1_n58), .A2(
        mul_y0y1_gf4_mul_1_1_n60), .ZN(mul_y0y1_gf4_mul_1_1_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_1_1_U5 ( .A(Y0xD[5]), .B(Y0xD[7]), .Z(
        mul_y0y1_gf4_mul_1_1_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_1_1_U4 ( .A(Y1xD[5]), .B(Y1xD[7]), .Z(
        mul_y0y1_gf4_mul_1_1_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_1_1_U3 ( .A1(mul_y0y1_gf4_mul_1_1_n54), .A2(
        mul_y0y1_gf4_mul_1_1_n53), .ZN(mul_y0y1_gf4_mul_1_1_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U2 ( .A(Y1xD[4]), .B(Y1xD[5]), .ZN(
        mul_y0y1_gf4_mul_1_1_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_1_U1 ( .A(Y0xD[4]), .B(Y0xD[5]), .ZN(
        mul_y0y1_gf4_mul_1_1_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U29 ( .A(mul_y0y1_gf4_mul_1_0_n77), .B(
        mul_y0y1_gf4_mul_1_0_n76), .ZN(mul_y0y1_Xi_mul_Yj_4__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_0_U28 ( .A1(Y1xD[7]), .A2(Y0xD[3]), .ZN(
        mul_y0y1_gf4_mul_1_0_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_1_0_U27 ( .A(mul_y0y1_gf4_mul_1_0_n75), .B(
        mul_y0y1_gf4_mul_1_0_n74), .Z(mul_y0y1_gf4_mul_1_0_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U26 ( .A(mul_y0y1_gf4_mul_1_0_n73), .B(
        mul_y0y1_gf4_mul_1_0_n72), .ZN(mul_y0y1_Xi_mul_Yj_4__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_0_U25 ( .A1(Y1xD[6]), .A2(Y0xD[2]), .ZN(
        mul_y0y1_gf4_mul_1_0_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_1_0_U24 ( .A(mul_y0y1_gf4_mul_1_0_n74), .B(
        mul_y0y1_gf4_mul_1_0_n71), .Z(mul_y0y1_gf4_mul_1_0_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_1_0_U23 ( .A1(mul_y0y1_gf4_mul_1_0_n70), .A2(
        mul_y0y1_gf4_mul_1_0_n69), .ZN(mul_y0y1_gf4_mul_1_0_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U22 ( .A(Y1xD[6]), .B(Y1xD[7]), .ZN(
        mul_y0y1_gf4_mul_1_0_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U21 ( .A(Y0xD[2]), .B(Y0xD[3]), .ZN(
        mul_y0y1_gf4_mul_1_0_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U20 ( .A(mul_y0y1_gf4_mul_1_0_n68), .B(
        mul_y0y1_gf4_mul_1_0_n67), .ZN(mul_y0y1_Xi_mul_Yj_4__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_0_U19 ( .A1(Y1xD[5]), .A2(Y0xD[1]), .ZN(
        mul_y0y1_gf4_mul_1_0_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_1_0_U18 ( .A(mul_y0y1_gf4_mul_1_0_n75), .B(
        mul_y0y1_gf4_mul_1_0_n66), .Z(mul_y0y1_gf4_mul_1_0_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U17 ( .A(mul_y0y1_gf4_mul_1_0_n65), .B(
        mul_y0y1_gf4_mul_1_0_n64), .ZN(mul_y0y1_gf4_mul_1_0_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_1_0_U16 ( .A1(mul_y0y1_gf4_mul_1_0_n63), .A2(
        mul_y0y1_gf4_mul_1_0_n62), .ZN(mul_y0y1_gf4_mul_1_0_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U15 ( .A(mul_y0y1_gf4_mul_1_0_n61), .B(
        mul_y0y1_gf4_mul_1_0_n60), .ZN(mul_y0y1_gf4_mul_1_0_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U14 ( .A(mul_y0y1_gf4_mul_1_0_n59), .B(
        mul_y0y1_gf4_mul_1_0_n58), .ZN(mul_y0y1_gf4_mul_1_0_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U13 ( .A(mul_y0y1_gf4_mul_1_0_n57), .B(
        mul_y0y1_gf4_mul_1_0_n56), .ZN(mul_y0y1_Xi_mul_Yj_4__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_1_0_U12 ( .A1(Y1xD[4]), .A2(Y0xD[0]), .ZN(
        mul_y0y1_gf4_mul_1_0_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_1_0_U11 ( .A(mul_y0y1_gf4_mul_1_0_n66), .B(
        mul_y0y1_gf4_mul_1_0_n71), .Z(mul_y0y1_gf4_mul_1_0_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U10 ( .A(mul_y0y1_gf4_mul_1_0_n55), .B(
        mul_y0y1_gf4_mul_1_0_n65), .ZN(mul_y0y1_gf4_mul_1_0_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_1_0_U9 ( .A1(mul_y0y1_gf4_mul_1_0_n61), .A2(
        mul_y0y1_gf4_mul_1_0_n59), .ZN(mul_y0y1_gf4_mul_1_0_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U8 ( .A(Y1xD[4]), .B(Y1xD[6]), .ZN(
        mul_y0y1_gf4_mul_1_0_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U7 ( .A(Y0xD[0]), .B(Y0xD[2]), .ZN(
        mul_y0y1_gf4_mul_1_0_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_1_0_U6 ( .A1(mul_y0y1_gf4_mul_1_0_n58), .A2(
        mul_y0y1_gf4_mul_1_0_n60), .ZN(mul_y0y1_gf4_mul_1_0_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_1_0_U5 ( .A(Y0xD[1]), .B(Y0xD[3]), .Z(
        mul_y0y1_gf4_mul_1_0_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_1_0_U4 ( .A(Y1xD[5]), .B(Y1xD[7]), .Z(
        mul_y0y1_gf4_mul_1_0_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_1_0_U3 ( .A1(mul_y0y1_gf4_mul_1_0_n54), .A2(
        mul_y0y1_gf4_mul_1_0_n53), .ZN(mul_y0y1_gf4_mul_1_0_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U2 ( .A(Y1xD[4]), .B(Y1xD[5]), .ZN(
        mul_y0y1_gf4_mul_1_0_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_1_0_U1 ( .A(Y0xD[0]), .B(Y0xD[1]), .ZN(
        mul_y0y1_gf4_mul_1_0_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_3_U29 ( .A(mul_y0y1_gf4_mul_0_3_n77), .B(
        mul_y0y1_gf4_mul_0_3_n76), .ZN(mul_y0y1_Xi_mul_Yj_3__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_3_U28 ( .A1(Y1xD[3]), .A2(Y0xD[15]), .ZN(
        mul_y0y1_gf4_mul_0_3_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_0_3_U27 ( .A(mul_y0y1_gf4_mul_0_3_n75), .B(
        mul_y0y1_gf4_mul_0_3_n74), .Z(mul_y0y1_gf4_mul_0_3_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_3_U26 ( .A(mul_y0y1_gf4_mul_0_3_n73), .B(
        mul_y0y1_gf4_mul_0_3_n72), .ZN(mul_y0y1_Xi_mul_Yj_3__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_3_U25 ( .A1(Y1xD[2]), .A2(Y0xD[14]), .ZN(
        mul_y0y1_gf4_mul_0_3_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_0_3_U24 ( .A(mul_y0y1_gf4_mul_0_3_n74), .B(
        mul_y0y1_gf4_mul_0_3_n71), .Z(mul_y0y1_gf4_mul_0_3_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_0_3_U23 ( .A1(mul_y0y1_gf4_mul_0_3_n70), .A2(
        mul_y0y1_gf4_mul_0_3_n69), .ZN(mul_y0y1_gf4_mul_0_3_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_3_U22 ( .A(Y1xD[2]), .B(Y1xD[3]), .ZN(
        mul_y0y1_gf4_mul_0_3_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_3_U21 ( .A(Y0xD[14]), .B(Y0xD[15]), .ZN(
        mul_y0y1_gf4_mul_0_3_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_3_U20 ( .A(mul_y0y1_gf4_mul_0_3_n68), .B(
        mul_y0y1_gf4_mul_0_3_n67), .ZN(mul_y0y1_Xi_mul_Yj_3__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_3_U19 ( .A1(Y1xD[1]), .A2(Y0xD[13]), .ZN(
        mul_y0y1_gf4_mul_0_3_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_0_3_U18 ( .A(mul_y0y1_gf4_mul_0_3_n75), .B(
        mul_y0y1_gf4_mul_0_3_n66), .Z(mul_y0y1_gf4_mul_0_3_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_3_U17 ( .A(mul_y0y1_gf4_mul_0_3_n65), .B(
        mul_y0y1_gf4_mul_0_3_n64), .ZN(mul_y0y1_gf4_mul_0_3_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_0_3_U16 ( .A1(mul_y0y1_gf4_mul_0_3_n63), .A2(
        mul_y0y1_gf4_mul_0_3_n62), .ZN(mul_y0y1_gf4_mul_0_3_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_3_U15 ( .A(mul_y0y1_gf4_mul_0_3_n61), .B(
        mul_y0y1_gf4_mul_0_3_n60), .ZN(mul_y0y1_gf4_mul_0_3_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_3_U14 ( .A(mul_y0y1_gf4_mul_0_3_n59), .B(
        mul_y0y1_gf4_mul_0_3_n58), .ZN(mul_y0y1_gf4_mul_0_3_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_3_U13 ( .A(mul_y0y1_gf4_mul_0_3_n57), .B(
        mul_y0y1_gf4_mul_0_3_n56), .ZN(mul_y0y1_Xi_mul_Yj_3__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_3_U12 ( .A1(Y1xD[0]), .A2(Y0xD[12]), .ZN(
        mul_y0y1_gf4_mul_0_3_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_0_3_U11 ( .A(mul_y0y1_gf4_mul_0_3_n66), .B(
        mul_y0y1_gf4_mul_0_3_n71), .Z(mul_y0y1_gf4_mul_0_3_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_3_U10 ( .A(mul_y0y1_gf4_mul_0_3_n55), .B(
        mul_y0y1_gf4_mul_0_3_n65), .ZN(mul_y0y1_gf4_mul_0_3_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_0_3_U9 ( .A1(mul_y0y1_gf4_mul_0_3_n61), .A2(
        mul_y0y1_gf4_mul_0_3_n59), .ZN(mul_y0y1_gf4_mul_0_3_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_3_U8 ( .A(Y1xD[0]), .B(Y1xD[2]), .ZN(
        mul_y0y1_gf4_mul_0_3_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_3_U7 ( .A(Y0xD[12]), .B(Y0xD[14]), .ZN(
        mul_y0y1_gf4_mul_0_3_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_0_3_U6 ( .A1(mul_y0y1_gf4_mul_0_3_n58), .A2(
        mul_y0y1_gf4_mul_0_3_n60), .ZN(mul_y0y1_gf4_mul_0_3_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_0_3_U5 ( .A(Y0xD[13]), .B(Y0xD[15]), .Z(
        mul_y0y1_gf4_mul_0_3_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_0_3_U4 ( .A(Y1xD[1]), .B(Y1xD[3]), .Z(
        mul_y0y1_gf4_mul_0_3_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_0_3_U3 ( .A1(mul_y0y1_gf4_mul_0_3_n54), .A2(
        mul_y0y1_gf4_mul_0_3_n53), .ZN(mul_y0y1_gf4_mul_0_3_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_3_U2 ( .A(Y1xD[0]), .B(Y1xD[1]), .ZN(
        mul_y0y1_gf4_mul_0_3_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_3_U1 ( .A(Y0xD[12]), .B(Y0xD[13]), .ZN(
        mul_y0y1_gf4_mul_0_3_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U29 ( .A(mul_y0y1_gf4_mul_0_2_n77), .B(
        mul_y0y1_gf4_mul_0_2_n76), .ZN(mul_y0y1_Xi_mul_Yj_2__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_2_U28 ( .A1(Y1xD[3]), .A2(Y0xD[11]), .ZN(
        mul_y0y1_gf4_mul_0_2_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_0_2_U27 ( .A(mul_y0y1_gf4_mul_0_2_n75), .B(
        mul_y0y1_gf4_mul_0_2_n74), .Z(mul_y0y1_gf4_mul_0_2_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U26 ( .A(mul_y0y1_gf4_mul_0_2_n73), .B(
        mul_y0y1_gf4_mul_0_2_n72), .ZN(mul_y0y1_Xi_mul_Yj_2__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_2_U25 ( .A1(Y1xD[2]), .A2(Y0xD[10]), .ZN(
        mul_y0y1_gf4_mul_0_2_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_0_2_U24 ( .A(mul_y0y1_gf4_mul_0_2_n74), .B(
        mul_y0y1_gf4_mul_0_2_n71), .Z(mul_y0y1_gf4_mul_0_2_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_0_2_U23 ( .A1(mul_y0y1_gf4_mul_0_2_n70), .A2(
        mul_y0y1_gf4_mul_0_2_n69), .ZN(mul_y0y1_gf4_mul_0_2_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U22 ( .A(Y1xD[2]), .B(Y1xD[3]), .ZN(
        mul_y0y1_gf4_mul_0_2_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U21 ( .A(Y0xD[10]), .B(Y0xD[11]), .ZN(
        mul_y0y1_gf4_mul_0_2_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U20 ( .A(mul_y0y1_gf4_mul_0_2_n68), .B(
        mul_y0y1_gf4_mul_0_2_n67), .ZN(mul_y0y1_Xi_mul_Yj_2__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_2_U19 ( .A1(Y1xD[1]), .A2(Y0xD[9]), .ZN(
        mul_y0y1_gf4_mul_0_2_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_0_2_U18 ( .A(mul_y0y1_gf4_mul_0_2_n75), .B(
        mul_y0y1_gf4_mul_0_2_n66), .Z(mul_y0y1_gf4_mul_0_2_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U17 ( .A(mul_y0y1_gf4_mul_0_2_n65), .B(
        mul_y0y1_gf4_mul_0_2_n64), .ZN(mul_y0y1_gf4_mul_0_2_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_0_2_U16 ( .A1(mul_y0y1_gf4_mul_0_2_n63), .A2(
        mul_y0y1_gf4_mul_0_2_n62), .ZN(mul_y0y1_gf4_mul_0_2_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U15 ( .A(mul_y0y1_gf4_mul_0_2_n61), .B(
        mul_y0y1_gf4_mul_0_2_n60), .ZN(mul_y0y1_gf4_mul_0_2_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U14 ( .A(mul_y0y1_gf4_mul_0_2_n59), .B(
        mul_y0y1_gf4_mul_0_2_n58), .ZN(mul_y0y1_gf4_mul_0_2_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U13 ( .A(mul_y0y1_gf4_mul_0_2_n57), .B(
        mul_y0y1_gf4_mul_0_2_n56), .ZN(mul_y0y1_Xi_mul_Yj_2__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_2_U12 ( .A1(Y1xD[0]), .A2(Y0xD[8]), .ZN(
        mul_y0y1_gf4_mul_0_2_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_0_2_U11 ( .A(mul_y0y1_gf4_mul_0_2_n66), .B(
        mul_y0y1_gf4_mul_0_2_n71), .Z(mul_y0y1_gf4_mul_0_2_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U10 ( .A(mul_y0y1_gf4_mul_0_2_n55), .B(
        mul_y0y1_gf4_mul_0_2_n65), .ZN(mul_y0y1_gf4_mul_0_2_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_0_2_U9 ( .A1(mul_y0y1_gf4_mul_0_2_n61), .A2(
        mul_y0y1_gf4_mul_0_2_n59), .ZN(mul_y0y1_gf4_mul_0_2_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U8 ( .A(Y1xD[0]), .B(Y1xD[2]), .ZN(
        mul_y0y1_gf4_mul_0_2_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U7 ( .A(Y0xD[8]), .B(Y0xD[10]), .ZN(
        mul_y0y1_gf4_mul_0_2_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_0_2_U6 ( .A1(mul_y0y1_gf4_mul_0_2_n58), .A2(
        mul_y0y1_gf4_mul_0_2_n60), .ZN(mul_y0y1_gf4_mul_0_2_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_0_2_U5 ( .A(Y0xD[9]), .B(Y0xD[11]), .Z(
        mul_y0y1_gf4_mul_0_2_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_0_2_U4 ( .A(Y1xD[1]), .B(Y1xD[3]), .Z(
        mul_y0y1_gf4_mul_0_2_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_0_2_U3 ( .A1(mul_y0y1_gf4_mul_0_2_n54), .A2(
        mul_y0y1_gf4_mul_0_2_n53), .ZN(mul_y0y1_gf4_mul_0_2_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U2 ( .A(Y1xD[0]), .B(Y1xD[1]), .ZN(
        mul_y0y1_gf4_mul_0_2_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_2_U1 ( .A(Y0xD[8]), .B(Y0xD[9]), .ZN(
        mul_y0y1_gf4_mul_0_2_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U29 ( .A(mul_y0y1_gf4_mul_0_1_n77), .B(
        mul_y0y1_gf4_mul_0_1_n76), .ZN(mul_y0y1_Xi_mul_Yj_1__3_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_1_U28 ( .A1(Y1xD[3]), .A2(Y0xD[7]), .ZN(
        mul_y0y1_gf4_mul_0_1_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_0_1_U27 ( .A(mul_y0y1_gf4_mul_0_1_n75), .B(
        mul_y0y1_gf4_mul_0_1_n74), .Z(mul_y0y1_gf4_mul_0_1_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U26 ( .A(mul_y0y1_gf4_mul_0_1_n73), .B(
        mul_y0y1_gf4_mul_0_1_n72), .ZN(mul_y0y1_Xi_mul_Yj_1__2_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_1_U25 ( .A1(Y1xD[2]), .A2(Y0xD[6]), .ZN(
        mul_y0y1_gf4_mul_0_1_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_0_1_U24 ( .A(mul_y0y1_gf4_mul_0_1_n74), .B(
        mul_y0y1_gf4_mul_0_1_n71), .Z(mul_y0y1_gf4_mul_0_1_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_0_1_U23 ( .A1(mul_y0y1_gf4_mul_0_1_n70), .A2(
        mul_y0y1_gf4_mul_0_1_n69), .ZN(mul_y0y1_gf4_mul_0_1_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U22 ( .A(Y1xD[2]), .B(Y1xD[3]), .ZN(
        mul_y0y1_gf4_mul_0_1_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U21 ( .A(Y0xD[6]), .B(Y0xD[7]), .ZN(
        mul_y0y1_gf4_mul_0_1_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U20 ( .A(mul_y0y1_gf4_mul_0_1_n68), .B(
        mul_y0y1_gf4_mul_0_1_n67), .ZN(mul_y0y1_Xi_mul_Yj_1__1_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_1_U19 ( .A1(Y1xD[1]), .A2(Y0xD[5]), .ZN(
        mul_y0y1_gf4_mul_0_1_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_0_1_U18 ( .A(mul_y0y1_gf4_mul_0_1_n75), .B(
        mul_y0y1_gf4_mul_0_1_n66), .Z(mul_y0y1_gf4_mul_0_1_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U17 ( .A(mul_y0y1_gf4_mul_0_1_n65), .B(
        mul_y0y1_gf4_mul_0_1_n64), .ZN(mul_y0y1_gf4_mul_0_1_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_0_1_U16 ( .A1(mul_y0y1_gf4_mul_0_1_n63), .A2(
        mul_y0y1_gf4_mul_0_1_n62), .ZN(mul_y0y1_gf4_mul_0_1_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U15 ( .A(mul_y0y1_gf4_mul_0_1_n61), .B(
        mul_y0y1_gf4_mul_0_1_n60), .ZN(mul_y0y1_gf4_mul_0_1_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U14 ( .A(mul_y0y1_gf4_mul_0_1_n59), .B(
        mul_y0y1_gf4_mul_0_1_n58), .ZN(mul_y0y1_gf4_mul_0_1_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U13 ( .A(mul_y0y1_gf4_mul_0_1_n57), .B(
        mul_y0y1_gf4_mul_0_1_n56), .ZN(mul_y0y1_Xi_mul_Yj_1__0_) );
  NAND2_X1 mul_y0y1_gf4_mul_0_1_U12 ( .A1(Y1xD[0]), .A2(Y0xD[4]), .ZN(
        mul_y0y1_gf4_mul_0_1_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_0_1_U11 ( .A(mul_y0y1_gf4_mul_0_1_n66), .B(
        mul_y0y1_gf4_mul_0_1_n71), .Z(mul_y0y1_gf4_mul_0_1_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U10 ( .A(mul_y0y1_gf4_mul_0_1_n55), .B(
        mul_y0y1_gf4_mul_0_1_n65), .ZN(mul_y0y1_gf4_mul_0_1_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_0_1_U9 ( .A1(mul_y0y1_gf4_mul_0_1_n61), .A2(
        mul_y0y1_gf4_mul_0_1_n59), .ZN(mul_y0y1_gf4_mul_0_1_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U8 ( .A(Y1xD[0]), .B(Y1xD[2]), .ZN(
        mul_y0y1_gf4_mul_0_1_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U7 ( .A(Y0xD[4]), .B(Y0xD[6]), .ZN(
        mul_y0y1_gf4_mul_0_1_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_0_1_U6 ( .A1(mul_y0y1_gf4_mul_0_1_n58), .A2(
        mul_y0y1_gf4_mul_0_1_n60), .ZN(mul_y0y1_gf4_mul_0_1_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_0_1_U5 ( .A(Y0xD[5]), .B(Y0xD[7]), .Z(
        mul_y0y1_gf4_mul_0_1_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_0_1_U4 ( .A(Y1xD[1]), .B(Y1xD[3]), .Z(
        mul_y0y1_gf4_mul_0_1_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_0_1_U3 ( .A1(mul_y0y1_gf4_mul_0_1_n54), .A2(
        mul_y0y1_gf4_mul_0_1_n53), .ZN(mul_y0y1_gf4_mul_0_1_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U2 ( .A(Y1xD[0]), .B(Y1xD[1]), .ZN(
        mul_y0y1_gf4_mul_0_1_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_1_U1 ( .A(Y0xD[4]), .B(Y0xD[5]), .ZN(
        mul_y0y1_gf4_mul_0_1_n54) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U29 ( .A(mul_y0y1_gf4_mul_0_0_n77), .B(
        mul_y0y1_gf4_mul_0_0_n76), .ZN(mul_y0y1_FFxDN[3]) );
  NAND2_X1 mul_y0y1_gf4_mul_0_0_U28 ( .A1(Y1xD[3]), .A2(Y0xD[3]), .ZN(
        mul_y0y1_gf4_mul_0_0_n76) );
  XOR2_X1 mul_y0y1_gf4_mul_0_0_U27 ( .A(mul_y0y1_gf4_mul_0_0_n75), .B(
        mul_y0y1_gf4_mul_0_0_n74), .Z(mul_y0y1_gf4_mul_0_0_n77) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U26 ( .A(mul_y0y1_gf4_mul_0_0_n73), .B(
        mul_y0y1_gf4_mul_0_0_n72), .ZN(mul_y0y1_FFxDN[2]) );
  NAND2_X1 mul_y0y1_gf4_mul_0_0_U25 ( .A1(Y1xD[2]), .A2(Y0xD[2]), .ZN(
        mul_y0y1_gf4_mul_0_0_n72) );
  XOR2_X1 mul_y0y1_gf4_mul_0_0_U24 ( .A(mul_y0y1_gf4_mul_0_0_n74), .B(
        mul_y0y1_gf4_mul_0_0_n71), .Z(mul_y0y1_gf4_mul_0_0_n73) );
  NOR2_X1 mul_y0y1_gf4_mul_0_0_U23 ( .A1(mul_y0y1_gf4_mul_0_0_n70), .A2(
        mul_y0y1_gf4_mul_0_0_n69), .ZN(mul_y0y1_gf4_mul_0_0_n74) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U22 ( .A(Y1xD[2]), .B(Y1xD[3]), .ZN(
        mul_y0y1_gf4_mul_0_0_n69) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U21 ( .A(Y0xD[2]), .B(Y0xD[3]), .ZN(
        mul_y0y1_gf4_mul_0_0_n70) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U20 ( .A(mul_y0y1_gf4_mul_0_0_n68), .B(
        mul_y0y1_gf4_mul_0_0_n67), .ZN(mul_y0y1_FFxDN[1]) );
  NAND2_X1 mul_y0y1_gf4_mul_0_0_U19 ( .A1(Y1xD[1]), .A2(Y0xD[1]), .ZN(
        mul_y0y1_gf4_mul_0_0_n67) );
  XOR2_X1 mul_y0y1_gf4_mul_0_0_U18 ( .A(mul_y0y1_gf4_mul_0_0_n75), .B(
        mul_y0y1_gf4_mul_0_0_n66), .Z(mul_y0y1_gf4_mul_0_0_n68) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U17 ( .A(mul_y0y1_gf4_mul_0_0_n65), .B(
        mul_y0y1_gf4_mul_0_0_n64), .ZN(mul_y0y1_gf4_mul_0_0_n75) );
  NAND2_X1 mul_y0y1_gf4_mul_0_0_U16 ( .A1(mul_y0y1_gf4_mul_0_0_n63), .A2(
        mul_y0y1_gf4_mul_0_0_n62), .ZN(mul_y0y1_gf4_mul_0_0_n64) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U15 ( .A(mul_y0y1_gf4_mul_0_0_n61), .B(
        mul_y0y1_gf4_mul_0_0_n60), .ZN(mul_y0y1_gf4_mul_0_0_n62) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U14 ( .A(mul_y0y1_gf4_mul_0_0_n59), .B(
        mul_y0y1_gf4_mul_0_0_n58), .ZN(mul_y0y1_gf4_mul_0_0_n63) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U13 ( .A(mul_y0y1_gf4_mul_0_0_n57), .B(
        mul_y0y1_gf4_mul_0_0_n56), .ZN(mul_y0y1_FFxDN[0]) );
  NAND2_X1 mul_y0y1_gf4_mul_0_0_U12 ( .A1(Y1xD[0]), .A2(Y0xD[0]), .ZN(
        mul_y0y1_gf4_mul_0_0_n56) );
  XOR2_X1 mul_y0y1_gf4_mul_0_0_U11 ( .A(mul_y0y1_gf4_mul_0_0_n66), .B(
        mul_y0y1_gf4_mul_0_0_n71), .Z(mul_y0y1_gf4_mul_0_0_n57) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U10 ( .A(mul_y0y1_gf4_mul_0_0_n55), .B(
        mul_y0y1_gf4_mul_0_0_n65), .ZN(mul_y0y1_gf4_mul_0_0_n71) );
  NOR2_X1 mul_y0y1_gf4_mul_0_0_U9 ( .A1(mul_y0y1_gf4_mul_0_0_n61), .A2(
        mul_y0y1_gf4_mul_0_0_n59), .ZN(mul_y0y1_gf4_mul_0_0_n65) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U8 ( .A(Y1xD[0]), .B(Y1xD[2]), .ZN(
        mul_y0y1_gf4_mul_0_0_n59) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U7 ( .A(Y0xD[0]), .B(Y0xD[2]), .ZN(
        mul_y0y1_gf4_mul_0_0_n61) );
  NAND2_X1 mul_y0y1_gf4_mul_0_0_U6 ( .A1(mul_y0y1_gf4_mul_0_0_n58), .A2(
        mul_y0y1_gf4_mul_0_0_n60), .ZN(mul_y0y1_gf4_mul_0_0_n55) );
  XOR2_X1 mul_y0y1_gf4_mul_0_0_U5 ( .A(Y0xD[1]), .B(Y0xD[3]), .Z(
        mul_y0y1_gf4_mul_0_0_n60) );
  XOR2_X1 mul_y0y1_gf4_mul_0_0_U4 ( .A(Y1xD[1]), .B(Y1xD[3]), .Z(
        mul_y0y1_gf4_mul_0_0_n58) );
  NOR2_X1 mul_y0y1_gf4_mul_0_0_U3 ( .A1(mul_y0y1_gf4_mul_0_0_n54), .A2(
        mul_y0y1_gf4_mul_0_0_n53), .ZN(mul_y0y1_gf4_mul_0_0_n66) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U2 ( .A(Y1xD[0]), .B(Y1xD[1]), .ZN(
        mul_y0y1_gf4_mul_0_0_n53) );
  XNOR2_X1 mul_y0y1_gf4_mul_0_0_U1 ( .A(Y0xD[0]), .B(Y0xD[1]), .ZN(
        mul_y0y1_gf4_mul_0_0_n54) );
  XNOR2_X1 inverter_gf24_U23 ( .A(inverter_gf24_n4), .B(InverterInxDP[14]), 
        .ZN(inverter_gf24_n13) );
  XNOR2_X1 inverter_gf24_U22 ( .A(inverter_gf24_d_3__0_), .B(InverterInxDP[12]), .ZN(inverter_gf24_n4) );
  XNOR2_X1 inverter_gf24_U21 ( .A(inverter_gf24_n3), .B(InverterInxDP[10]), 
        .ZN(inverter_gf24_n14) );
  XNOR2_X1 inverter_gf24_U20 ( .A(inverter_gf24_d_2__0_), .B(InverterInxDP[8]), 
        .ZN(inverter_gf24_n3) );
  XNOR2_X1 inverter_gf24_U19 ( .A(inverter_gf24_n2), .B(InverterInxDP[6]), 
        .ZN(inverter_gf24_n15) );
  XNOR2_X1 inverter_gf24_U18 ( .A(inverter_gf24_d_1__0_), .B(InverterInxDP[4]), 
        .ZN(inverter_gf24_n2) );
  XNOR2_X1 inverter_gf24_U17 ( .A(inverter_gf24_n1), .B(InverterInxDP[2]), 
        .ZN(inverter_gf24_n16) );
  XNOR2_X1 inverter_gf24_U16 ( .A(inverter_gf24_d_0__0_), .B(InverterInxDP[0]), 
        .ZN(inverter_gf24_n1) );
  XOR2_X1 inverter_gf24_U15 ( .A(InverterInxDP[13]), .B(InverterInxDP[15]), 
        .Z(inverter_gf24_d_3__0_) );
  XOR2_X1 inverter_gf24_U14 ( .A(InverterInxDP[9]), .B(InverterInxDP[11]), .Z(
        inverter_gf24_d_2__0_) );
  XOR2_X1 inverter_gf24_U13 ( .A(InverterInxDP[5]), .B(InverterInxDP[7]), .Z(
        inverter_gf24_d_1__0_) );
  XOR2_X1 inverter_gf24_U12 ( .A(InverterInxDP[1]), .B(InverterInxDP[3]), .Z(
        inverter_gf24_d_0__0_) );
  XNOR2_X1 inverter_gf24_U11 ( .A(inverter_gf24_AmulBxD[6]), .B(
        inverter_gf24_n5), .ZN(inverter_gf24_ExD[7]) );
  XNOR2_X1 inverter_gf24_U10 ( .A(inverter_gf24_AmulBxD[7]), .B(
        inverter_gf24_n6), .ZN(inverter_gf24_ExD[6]) );
  XNOR2_X1 inverter_gf24_U9 ( .A(inverter_gf24_AmulBxD[4]), .B(
        inverter_gf24_n7), .ZN(inverter_gf24_ExD[5]) );
  XNOR2_X1 inverter_gf24_U8 ( .A(inverter_gf24_AmulBxD[5]), .B(
        inverter_gf24_n8), .ZN(inverter_gf24_ExD[4]) );
  XNOR2_X1 inverter_gf24_U7 ( .A(inverter_gf24_AmulBxD[2]), .B(
        inverter_gf24_n9), .ZN(inverter_gf24_ExD[3]) );
  XNOR2_X1 inverter_gf24_U6 ( .A(inverter_gf24_AmulBxD[3]), .B(
        inverter_gf24_n10), .ZN(inverter_gf24_ExD[2]) );
  XNOR2_X1 inverter_gf24_U5 ( .A(inverter_gf24_AmulBxD[0]), .B(
        inverter_gf24_n11), .ZN(inverter_gf24_ExD[1]) );
  XNOR2_X1 inverter_gf24_U4 ( .A(inverter_gf24_AmulBxD[1]), .B(
        inverter_gf24_n12), .ZN(inverter_gf24_ExD[0]) );
  DFF_X1 inverter_gf24_CxDP_reg_0__0_ ( .D(inverter_gf24_n16), .CK(ClkxCI), 
        .Q(), .QN(inverter_gf24_n11) );
  DFF_X1 inverter_gf24_CxDP_reg_1__0_ ( .D(inverter_gf24_n15), .CK(ClkxCI), 
        .Q(), .QN(inverter_gf24_n9) );
  DFF_X1 inverter_gf24_CxDP_reg_2__0_ ( .D(inverter_gf24_n14), .CK(ClkxCI), 
        .Q(), .QN(inverter_gf24_n7) );
  DFF_X1 inverter_gf24_CxDP_reg_3__0_ ( .D(inverter_gf24_n13), .CK(ClkxCI), 
        .Q(), .QN(inverter_gf24_n5) );
  DFF_X1 inverter_gf24_CxDP_reg_0__1_ ( .D(inverter_gf24_d_0__0_), .CK(ClkxCI), 
        .Q(), .QN(inverter_gf24_n12) );
  DFF_X1 inverter_gf24_CxDP_reg_1__1_ ( .D(inverter_gf24_d_1__0_), .CK(ClkxCI), 
        .Q(), .QN(inverter_gf24_n10) );
  DFF_X1 inverter_gf24_CxDP_reg_2__1_ ( .D(inverter_gf24_d_2__0_), .CK(ClkxCI), 
        .Q(), .QN(inverter_gf24_n8) );
  DFF_X1 inverter_gf24_CxDP_reg_3__1_ ( .D(inverter_gf24_d_3__0_), .CK(ClkxCI), 
        .Q(), .QN(inverter_gf24_n6) );
  DFF_X1 inverter_gf24_ExDP_reg_0__0_ ( .D(inverter_gf24_ExD[0]), .CK(ClkxCI), 
        .Q(inverter_gf24_ExDP_0__0_), .QN() );
  DFF_X1 inverter_gf24_ExDP_reg_0__1_ ( .D(inverter_gf24_ExD[1]), .CK(ClkxCI), 
        .Q(inverter_gf24_ExDP_0__1_), .QN() );
  DFF_X1 inverter_gf24_ExDP_reg_1__0_ ( .D(inverter_gf24_ExD[2]), .CK(ClkxCI), 
        .Q(inverter_gf24_ExDP_1__0_), .QN() );
  DFF_X1 inverter_gf24_ExDP_reg_1__1_ ( .D(inverter_gf24_ExD[3]), .CK(ClkxCI), 
        .Q(inverter_gf24_ExDP_1__1_), .QN() );
  DFF_X1 inverter_gf24_ExDP_reg_2__0_ ( .D(inverter_gf24_ExD[4]), .CK(ClkxCI), 
        .Q(inverter_gf24_ExDP_2__0_), .QN() );
  DFF_X1 inverter_gf24_ExDP_reg_2__1_ ( .D(inverter_gf24_ExD[5]), .CK(ClkxCI), 
        .Q(inverter_gf24_ExDP_2__1_), .QN() );
  DFF_X1 inverter_gf24_ExDP_reg_3__0_ ( .D(inverter_gf24_ExD[6]), .CK(ClkxCI), 
        .Q(inverter_gf24_ExDP_3__0_), .QN() );
  DFF_X1 inverter_gf24_ExDP_reg_3__1_ ( .D(inverter_gf24_ExD[7]), .CK(ClkxCI), 
        .Q(inverter_gf24_ExDP_3__1_), .QN() );
  DFF_X1 inverter_gf24_BxDP_reg_0__0_ ( .D(InverterInxDP[0]), .CK(ClkxCI), .Q(
        inverter_gf24_BxDP[0]), .QN() );
  DFF_X1 inverter_gf24_BxDP_reg_1__0_ ( .D(InverterInxDP[4]), .CK(ClkxCI), .Q(
        inverter_gf24_BxDP[2]), .QN() );
  DFF_X1 inverter_gf24_BxDP_reg_2__0_ ( .D(InverterInxDP[8]), .CK(ClkxCI), .Q(
        inverter_gf24_BxDP[4]), .QN() );
  DFF_X1 inverter_gf24_BxDP_reg_3__0_ ( .D(InverterInxDP[12]), .CK(ClkxCI), 
        .Q(inverter_gf24_BxDP[6]), .QN() );
  DFF_X1 inverter_gf24_AxDP_reg_0__0_ ( .D(InverterInxDP[2]), .CK(ClkxCI), .Q(
        inverter_gf24_AxDP[0]), .QN() );
  DFF_X1 inverter_gf24_AxDP_reg_1__0_ ( .D(InverterInxDP[6]), .CK(ClkxCI), .Q(
        inverter_gf24_AxDP[2]), .QN() );
  DFF_X1 inverter_gf24_AxDP_reg_2__0_ ( .D(InverterInxDP[10]), .CK(ClkxCI), 
        .Q(inverter_gf24_AxDP[4]), .QN() );
  DFF_X1 inverter_gf24_AxDP_reg_3__0_ ( .D(InverterInxDP[14]), .CK(ClkxCI), 
        .Q(inverter_gf24_AxDP[6]), .QN() );
  DFF_X1 inverter_gf24_AxDP_reg_0__1_ ( .D(InverterInxDP[3]), .CK(ClkxCI), .Q(
        inverter_gf24_AxDP[1]), .QN() );
  DFF_X1 inverter_gf24_AxDP_reg_1__1_ ( .D(InverterInxDP[7]), .CK(ClkxCI), .Q(
        inverter_gf24_AxDP[3]), .QN() );
  DFF_X1 inverter_gf24_AxDP_reg_2__1_ ( .D(InverterInxDP[11]), .CK(ClkxCI), 
        .Q(inverter_gf24_AxDP[5]), .QN() );
  DFF_X1 inverter_gf24_AxDP_reg_3__1_ ( .D(InverterInxDP[15]), .CK(ClkxCI), 
        .Q(inverter_gf24_AxDP[7]), .QN() );
  DFF_X1 inverter_gf24_BxDP_reg_0__1_ ( .D(InverterInxDP[1]), .CK(ClkxCI), .Q(
        inverter_gf24_BxDP[1]), .QN() );
  DFF_X1 inverter_gf24_BxDP_reg_1__1_ ( .D(InverterInxDP[5]), .CK(ClkxCI), .Q(
        inverter_gf24_BxDP[3]), .QN() );
  DFF_X1 inverter_gf24_BxDP_reg_2__1_ ( .D(InverterInxDP[9]), .CK(ClkxCI), .Q(
        inverter_gf24_BxDP[5]), .QN() );
  DFF_X1 inverter_gf24_BxDP_reg_3__1_ ( .D(InverterInxDP[13]), .CK(ClkxCI), 
        .Q(inverter_gf24_BxDP[7]), .QN() );
  DFF_X1 inverter_gf24_pipelinedAxDP_reg_0__0_ ( .D(inverter_gf24_AxDP[0]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedAxDP[0]), .QN() );
  DFF_X1 inverter_gf24_pipelinedAxDP_reg_0__1_ ( .D(inverter_gf24_AxDP[1]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedAxDP[1]), .QN() );
  DFF_X1 inverter_gf24_pipelinedAxDP_reg_1__0_ ( .D(inverter_gf24_AxDP[2]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedAxDP[2]), .QN() );
  DFF_X1 inverter_gf24_pipelinedAxDP_reg_1__1_ ( .D(inverter_gf24_AxDP[3]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedAxDP[3]), .QN() );
  DFF_X1 inverter_gf24_pipelinedAxDP_reg_2__0_ ( .D(inverter_gf24_AxDP[4]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedAxDP[4]), .QN() );
  DFF_X1 inverter_gf24_pipelinedAxDP_reg_2__1_ ( .D(inverter_gf24_AxDP[5]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedAxDP[5]), .QN() );
  DFF_X1 inverter_gf24_pipelinedAxDP_reg_3__0_ ( .D(inverter_gf24_AxDP[6]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedAxDP[6]), .QN() );
  DFF_X1 inverter_gf24_pipelinedAxDP_reg_3__1_ ( .D(inverter_gf24_AxDP[7]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedAxDP[7]), .QN() );
  DFF_X1 inverter_gf24_pipelinedBxDP_reg_0__0_ ( .D(inverter_gf24_BxDP[0]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedBxDP[0]), .QN() );
  DFF_X1 inverter_gf24_pipelinedBxDP_reg_0__1_ ( .D(inverter_gf24_BxDP[1]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedBxDP[1]), .QN() );
  DFF_X1 inverter_gf24_pipelinedBxDP_reg_1__0_ ( .D(inverter_gf24_BxDP[2]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedBxDP[2]), .QN() );
  DFF_X1 inverter_gf24_pipelinedBxDP_reg_1__1_ ( .D(inverter_gf24_BxDP[3]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedBxDP[3]), .QN() );
  DFF_X1 inverter_gf24_pipelinedBxDP_reg_2__0_ ( .D(inverter_gf24_BxDP[4]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedBxDP[4]), .QN() );
  DFF_X1 inverter_gf24_pipelinedBxDP_reg_2__1_ ( .D(inverter_gf24_BxDP[5]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedBxDP[5]), .QN() );
  DFF_X1 inverter_gf24_pipelinedBxDP_reg_3__0_ ( .D(inverter_gf24_BxDP[6]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedBxDP[6]), .QN() );
  DFF_X1 inverter_gf24_pipelinedBxDP_reg_3__1_ ( .D(inverter_gf24_BxDP[7]), 
        .CK(ClkxCI), .Q(inverter_gf24_pipelinedBxDP[7]), .QN() );
  XNOR2_X1 inverter_gf24_a_mul_b_U50 ( .A(inverter_gf24_a_mul_b_n16), .B(
        inverter_gf24_a_mul_b_n15), .ZN(inverter_gf24_AmulBxD[7]) );
  XNOR2_X1 inverter_gf24_a_mul_b_U49 ( .A(inverter_gf24_a_mul_b_n18), .B(
        inverter_gf24_a_mul_b_n17), .ZN(inverter_gf24_a_mul_b_n15) );
  XOR2_X1 inverter_gf24_a_mul_b_U48 ( .A(inverter_gf24_a_mul_b_n20), .B(
        inverter_gf24_a_mul_b_n19), .Z(inverter_gf24_a_mul_b_n16) );
  XNOR2_X1 inverter_gf24_a_mul_b_U47 ( .A(inverter_gf24_a_mul_b_n14), .B(
        inverter_gf24_a_mul_b_n13), .ZN(inverter_gf24_AmulBxD[6]) );
  XNOR2_X1 inverter_gf24_a_mul_b_U46 ( .A(inverter_gf24_a_mul_b_n22), .B(
        inverter_gf24_a_mul_b_n21), .ZN(inverter_gf24_a_mul_b_n13) );
  XOR2_X1 inverter_gf24_a_mul_b_U45 ( .A(inverter_gf24_a_mul_b_n24), .B(
        inverter_gf24_a_mul_b_n23), .Z(inverter_gf24_a_mul_b_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_U44 ( .A(inverter_gf24_a_mul_b_n12), .B(
        inverter_gf24_a_mul_b_n11), .ZN(inverter_gf24_AmulBxD[5]) );
  XNOR2_X1 inverter_gf24_a_mul_b_U43 ( .A(inverter_gf24_a_mul_b_n26), .B(
        inverter_gf24_a_mul_b_n25), .ZN(inverter_gf24_a_mul_b_n11) );
  XOR2_X1 inverter_gf24_a_mul_b_U42 ( .A(inverter_gf24_a_mul_b_n28), .B(
        inverter_gf24_a_mul_b_n27), .Z(inverter_gf24_a_mul_b_n12) );
  XNOR2_X1 inverter_gf24_a_mul_b_U41 ( .A(inverter_gf24_a_mul_b_n10), .B(
        inverter_gf24_a_mul_b_n9), .ZN(inverter_gf24_AmulBxD[4]) );
  XNOR2_X1 inverter_gf24_a_mul_b_U40 ( .A(inverter_gf24_a_mul_b_n30), .B(
        inverter_gf24_a_mul_b_n29), .ZN(inverter_gf24_a_mul_b_n9) );
  XOR2_X1 inverter_gf24_a_mul_b_U39 ( .A(inverter_gf24_a_mul_b_n32), .B(
        inverter_gf24_a_mul_b_n31), .Z(inverter_gf24_a_mul_b_n10) );
  XNOR2_X1 inverter_gf24_a_mul_b_U38 ( .A(inverter_gf24_a_mul_b_n8), .B(
        inverter_gf24_a_mul_b_n7), .ZN(inverter_gf24_AmulBxD[3]) );
  XNOR2_X1 inverter_gf24_a_mul_b_U37 ( .A(inverter_gf24_a_mul_b_n34), .B(
        inverter_gf24_a_mul_b_n33), .ZN(inverter_gf24_a_mul_b_n7) );
  XOR2_X1 inverter_gf24_a_mul_b_U36 ( .A(inverter_gf24_a_mul_b_n36), .B(
        inverter_gf24_a_mul_b_n35), .Z(inverter_gf24_a_mul_b_n8) );
  XNOR2_X1 inverter_gf24_a_mul_b_U35 ( .A(inverter_gf24_a_mul_b_n6), .B(
        inverter_gf24_a_mul_b_n5), .ZN(inverter_gf24_AmulBxD[2]) );
  XNOR2_X1 inverter_gf24_a_mul_b_U34 ( .A(inverter_gf24_a_mul_b_n38), .B(
        inverter_gf24_a_mul_b_n37), .ZN(inverter_gf24_a_mul_b_n5) );
  XOR2_X1 inverter_gf24_a_mul_b_U33 ( .A(inverter_gf24_a_mul_b_n40), .B(
        inverter_gf24_a_mul_b_n39), .Z(inverter_gf24_a_mul_b_n6) );
  XNOR2_X1 inverter_gf24_a_mul_b_U32 ( .A(inverter_gf24_a_mul_b_n4), .B(
        inverter_gf24_a_mul_b_n3), .ZN(inverter_gf24_AmulBxD[1]) );
  XNOR2_X1 inverter_gf24_a_mul_b_U31 ( .A(inverter_gf24_a_mul_b_n42), .B(
        inverter_gf24_a_mul_b_n41), .ZN(inverter_gf24_a_mul_b_n3) );
  XOR2_X1 inverter_gf24_a_mul_b_U30 ( .A(inverter_gf24_a_mul_b_n44), .B(
        inverter_gf24_a_mul_b_n43), .Z(inverter_gf24_a_mul_b_n4) );
  XNOR2_X1 inverter_gf24_a_mul_b_U29 ( .A(inverter_gf24_a_mul_b_n2), .B(
        inverter_gf24_a_mul_b_n1), .ZN(inverter_gf24_AmulBxD[0]) );
  XNOR2_X1 inverter_gf24_a_mul_b_U28 ( .A(inverter_gf24_a_mul_b_n46), .B(
        inverter_gf24_a_mul_b_n45), .ZN(inverter_gf24_a_mul_b_n1) );
  XOR2_X1 inverter_gf24_a_mul_b_U27 ( .A(inverter_gf24_a_mul_b_n48), .B(
        inverter_gf24_a_mul_b_n47), .Z(inverter_gf24_a_mul_b_n2) );
  XOR2_X1 inverter_gf24_a_mul_b_U26 ( .A(Zinv1xDI[5]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_9__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[19]) );
  XOR2_X1 inverter_gf24_a_mul_b_U25 ( .A(Zinv1xDI[4]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_9__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[18]) );
  XOR2_X1 inverter_gf24_a_mul_b_U24 ( .A(Zinv1xDI[3]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_8__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[17]) );
  XOR2_X1 inverter_gf24_a_mul_b_U23 ( .A(Zinv1xDI[2]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_8__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[16]) );
  XOR2_X1 inverter_gf24_a_mul_b_U22 ( .A(Zinv1xDI[9]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_7__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[15]) );
  XOR2_X1 inverter_gf24_a_mul_b_U21 ( .A(Zinv1xDI[8]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_7__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[14]) );
  XOR2_X1 inverter_gf24_a_mul_b_U20 ( .A(Zinv1xDI[5]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_6__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[13]) );
  XOR2_X1 inverter_gf24_a_mul_b_U19 ( .A(Zinv1xDI[4]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_6__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[12]) );
  XOR2_X1 inverter_gf24_a_mul_b_U18 ( .A(Zinv1xDI[1]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_4__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[9]) );
  XOR2_X1 inverter_gf24_a_mul_b_U17 ( .A(Zinv1xDI[0]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_4__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[8]) );
  XOR2_X1 inverter_gf24_a_mul_b_U16 ( .A(Zinv1xDI[7]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_3__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[7]) );
  XOR2_X1 inverter_gf24_a_mul_b_U15 ( .A(Zinv1xDI[6]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_3__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[6]) );
  XOR2_X1 inverter_gf24_a_mul_b_U14 ( .A(Zinv1xDI[3]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_2__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[5]) );
  XOR2_X1 inverter_gf24_a_mul_b_U13 ( .A(Zinv1xDI[2]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_2__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[4]) );
  XOR2_X1 inverter_gf24_a_mul_b_U12 ( .A(Zinv1xDI[1]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_1__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[3]) );
  XOR2_X1 inverter_gf24_a_mul_b_U11 ( .A(Zinv1xDI[0]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_1__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[2]) );
  XOR2_X1 inverter_gf24_a_mul_b_U10 ( .A(Zinv1xDI[11]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_14__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[29]) );
  XOR2_X1 inverter_gf24_a_mul_b_U9 ( .A(Zinv1xDI[10]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_14__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[28]) );
  XOR2_X1 inverter_gf24_a_mul_b_U8 ( .A(Zinv1xDI[9]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_13__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[27]) );
  XOR2_X1 inverter_gf24_a_mul_b_U7 ( .A(Zinv1xDI[8]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_13__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[26]) );
  XOR2_X1 inverter_gf24_a_mul_b_U6 ( .A(Zinv1xDI[7]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_12__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[25]) );
  XOR2_X1 inverter_gf24_a_mul_b_U5 ( .A(Zinv1xDI[6]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_12__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[24]) );
  XOR2_X1 inverter_gf24_a_mul_b_U4 ( .A(Zinv1xDI[11]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_11__1_), .Z(
        inverter_gf24_a_mul_b_FFxDN[23]) );
  XOR2_X1 inverter_gf24_a_mul_b_U3 ( .A(Zinv1xDI[10]), .B(
        inverter_gf24_a_mul_b_Xi_mul_Yj_11__0_), .Z(
        inverter_gf24_a_mul_b_FFxDN[22]) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_1__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[2]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n48) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_1__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[3]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n44) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_2__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[4]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n45) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_2__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[5]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n41) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_3__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[6]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n46) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_3__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[7]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n42) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_4__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[8]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n39) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_4__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[9]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n35) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_6__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[12]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n37) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_6__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[13]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n33) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_7__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[14]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n38) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_7__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[15]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n34) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_8__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[16]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n29) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_8__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[17]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n25) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_9__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[18]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n30) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_9__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[19]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n26) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_11__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[22]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n32) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_11__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[23]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n28) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_12__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[24]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n23) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_12__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[25]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n19) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_13__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[26]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n24) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_13__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[27]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n20) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_14__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[28]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n21) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_14__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[29]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n17) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_0__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[0]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n47) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_5__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[10]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n40) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_10__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[20]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n31) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_15__0_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[30]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n22) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_0__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[1]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n43) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_5__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[11]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n36) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_10__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[21]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n27) );
  DFF_X1 inverter_gf24_a_mul_b_FFxDP_reg_15__1_ ( .D(
        inverter_gf24_a_mul_b_FFxDN[31]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_b_n18) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_3_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_3_3_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_3_3_n14), .ZN(
        inverter_gf24_a_mul_b_FFxDN[31]) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_3_3_U6 ( .A1(InverterInxDP[15]), .A2(
        InverterInxDP[13]), .ZN(inverter_gf24_a_mul_b_gf2_mul_3_3_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_3_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_3_3_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_3_3_n14), .ZN(
        inverter_gf24_a_mul_b_FFxDN[30]) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_3_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_3_3_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_3_3_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_3_3_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_3_U3 ( .A(InverterInxDP[15]), .B(
        InverterInxDP[14]), .ZN(inverter_gf24_a_mul_b_gf2_mul_3_3_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_3_U2 ( .A(InverterInxDP[13]), .B(
        InverterInxDP[12]), .ZN(inverter_gf24_a_mul_b_gf2_mul_3_3_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_3_3_U1 ( .A1(InverterInxDP[14]), .A2(
        InverterInxDP[12]), .ZN(inverter_gf24_a_mul_b_gf2_mul_3_3_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_2_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_3_2_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_3_2_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_14__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_3_2_U6 ( .A1(InverterInxDP[15]), .A2(
        InverterInxDP[9]), .ZN(inverter_gf24_a_mul_b_gf2_mul_3_2_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_2_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_3_2_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_3_2_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_14__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_2_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_3_2_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_3_2_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_3_2_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_2_U3 ( .A(InverterInxDP[15]), .B(
        InverterInxDP[14]), .ZN(inverter_gf24_a_mul_b_gf2_mul_3_2_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_2_U2 ( .A(InverterInxDP[9]), .B(
        InverterInxDP[8]), .ZN(inverter_gf24_a_mul_b_gf2_mul_3_2_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_3_2_U1 ( .A1(InverterInxDP[14]), .A2(
        InverterInxDP[8]), .ZN(inverter_gf24_a_mul_b_gf2_mul_3_2_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_1_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_3_1_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_3_1_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_13__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_3_1_U6 ( .A1(InverterInxDP[15]), .A2(
        InverterInxDP[5]), .ZN(inverter_gf24_a_mul_b_gf2_mul_3_1_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_1_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_3_1_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_3_1_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_13__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_1_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_3_1_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_3_1_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_3_1_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_1_U3 ( .A(InverterInxDP[15]), .B(
        InverterInxDP[14]), .ZN(inverter_gf24_a_mul_b_gf2_mul_3_1_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_1_U2 ( .A(InverterInxDP[5]), .B(
        InverterInxDP[4]), .ZN(inverter_gf24_a_mul_b_gf2_mul_3_1_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_3_1_U1 ( .A1(InverterInxDP[14]), .A2(
        InverterInxDP[4]), .ZN(inverter_gf24_a_mul_b_gf2_mul_3_1_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_0_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_3_0_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_3_0_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_12__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_3_0_U6 ( .A1(InverterInxDP[15]), .A2(
        InverterInxDP[1]), .ZN(inverter_gf24_a_mul_b_gf2_mul_3_0_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_0_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_3_0_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_3_0_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_12__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_0_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_3_0_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_3_0_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_3_0_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_0_U3 ( .A(InverterInxDP[15]), .B(
        InverterInxDP[14]), .ZN(inverter_gf24_a_mul_b_gf2_mul_3_0_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_3_0_U2 ( .A(InverterInxDP[1]), .B(
        InverterInxDP[0]), .ZN(inverter_gf24_a_mul_b_gf2_mul_3_0_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_3_0_U1 ( .A1(InverterInxDP[14]), .A2(
        InverterInxDP[0]), .ZN(inverter_gf24_a_mul_b_gf2_mul_3_0_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_3_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_2_3_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_2_3_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_11__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_2_3_U6 ( .A1(InverterInxDP[11]), .A2(
        InverterInxDP[13]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_3_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_3_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_2_3_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_2_3_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_11__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_3_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_2_3_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_2_3_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_2_3_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_3_U3 ( .A(InverterInxDP[11]), .B(
        InverterInxDP[10]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_3_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_3_U2 ( .A(InverterInxDP[13]), .B(
        InverterInxDP[12]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_3_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_2_3_U1 ( .A1(InverterInxDP[10]), .A2(
        InverterInxDP[12]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_3_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_2_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_2_2_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_2_2_n14), .ZN(
        inverter_gf24_a_mul_b_FFxDN[21]) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_2_2_U6 ( .A1(InverterInxDP[11]), .A2(
        InverterInxDP[9]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_2_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_2_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_2_2_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_2_2_n14), .ZN(
        inverter_gf24_a_mul_b_FFxDN[20]) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_2_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_2_2_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_2_2_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_2_2_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_2_U3 ( .A(InverterInxDP[11]), .B(
        InverterInxDP[10]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_2_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_2_U2 ( .A(InverterInxDP[9]), .B(
        InverterInxDP[8]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_2_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_2_2_U1 ( .A1(InverterInxDP[10]), .A2(
        InverterInxDP[8]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_2_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_1_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_2_1_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_2_1_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_9__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_2_1_U6 ( .A1(InverterInxDP[11]), .A2(
        InverterInxDP[5]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_1_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_1_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_2_1_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_2_1_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_9__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_1_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_2_1_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_2_1_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_2_1_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_1_U3 ( .A(InverterInxDP[11]), .B(
        InverterInxDP[10]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_1_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_1_U2 ( .A(InverterInxDP[5]), .B(
        InverterInxDP[4]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_1_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_2_1_U1 ( .A1(InverterInxDP[10]), .A2(
        InverterInxDP[4]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_1_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_0_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_2_0_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_2_0_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_8__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_2_0_U6 ( .A1(InverterInxDP[11]), .A2(
        InverterInxDP[1]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_0_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_0_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_2_0_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_2_0_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_8__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_0_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_2_0_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_2_0_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_2_0_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_0_U3 ( .A(InverterInxDP[11]), .B(
        InverterInxDP[10]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_0_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_2_0_U2 ( .A(InverterInxDP[1]), .B(
        InverterInxDP[0]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_0_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_2_0_U1 ( .A1(InverterInxDP[10]), .A2(
        InverterInxDP[0]), .ZN(inverter_gf24_a_mul_b_gf2_mul_2_0_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_3_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_1_3_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_1_3_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_7__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_1_3_U6 ( .A1(InverterInxDP[7]), .A2(
        InverterInxDP[13]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_3_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_3_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_1_3_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_1_3_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_7__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_3_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_1_3_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_1_3_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_1_3_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_3_U3 ( .A(InverterInxDP[7]), .B(
        InverterInxDP[6]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_3_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_3_U2 ( .A(InverterInxDP[13]), .B(
        InverterInxDP[12]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_3_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_1_3_U1 ( .A1(InverterInxDP[6]), .A2(
        InverterInxDP[12]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_3_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_2_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_1_2_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_1_2_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_6__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_1_2_U6 ( .A1(InverterInxDP[7]), .A2(
        InverterInxDP[9]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_2_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_2_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_1_2_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_1_2_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_6__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_2_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_1_2_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_1_2_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_1_2_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_2_U3 ( .A(InverterInxDP[7]), .B(
        InverterInxDP[6]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_2_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_2_U2 ( .A(InverterInxDP[9]), .B(
        InverterInxDP[8]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_2_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_1_2_U1 ( .A1(InverterInxDP[6]), .A2(
        InverterInxDP[8]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_2_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_1_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_1_1_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_1_1_n14), .ZN(
        inverter_gf24_a_mul_b_FFxDN[11]) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_1_1_U6 ( .A1(InverterInxDP[7]), .A2(
        InverterInxDP[5]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_1_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_1_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_1_1_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_1_1_n14), .ZN(
        inverter_gf24_a_mul_b_FFxDN[10]) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_1_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_1_1_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_1_1_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_1_1_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_1_U3 ( .A(InverterInxDP[7]), .B(
        InverterInxDP[6]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_1_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_1_U2 ( .A(InverterInxDP[5]), .B(
        InverterInxDP[4]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_1_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_1_1_U1 ( .A1(InverterInxDP[6]), .A2(
        InverterInxDP[4]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_1_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_0_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_1_0_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_1_0_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_4__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_1_0_U6 ( .A1(InverterInxDP[7]), .A2(
        InverterInxDP[1]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_0_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_0_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_1_0_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_1_0_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_4__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_0_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_1_0_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_1_0_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_1_0_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_0_U3 ( .A(InverterInxDP[7]), .B(
        InverterInxDP[6]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_0_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_1_0_U2 ( .A(InverterInxDP[1]), .B(
        InverterInxDP[0]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_0_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_1_0_U1 ( .A1(InverterInxDP[6]), .A2(
        InverterInxDP[0]), .ZN(inverter_gf24_a_mul_b_gf2_mul_1_0_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_3_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_0_3_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_0_3_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_3__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_0_3_U6 ( .A1(InverterInxDP[3]), .A2(
        InverterInxDP[13]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_3_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_3_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_0_3_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_0_3_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_3__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_3_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_0_3_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_0_3_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_0_3_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_3_U3 ( .A(InverterInxDP[3]), .B(
        InverterInxDP[2]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_3_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_3_U2 ( .A(InverterInxDP[13]), .B(
        InverterInxDP[12]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_3_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_0_3_U1 ( .A1(InverterInxDP[2]), .A2(
        InverterInxDP[12]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_3_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_2_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_0_2_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_0_2_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_2__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_0_2_U6 ( .A1(InverterInxDP[3]), .A2(
        InverterInxDP[9]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_2_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_2_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_0_2_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_0_2_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_2__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_2_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_0_2_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_0_2_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_0_2_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_2_U3 ( .A(InverterInxDP[3]), .B(
        InverterInxDP[2]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_2_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_2_U2 ( .A(InverterInxDP[9]), .B(
        InverterInxDP[8]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_2_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_0_2_U1 ( .A1(InverterInxDP[2]), .A2(
        InverterInxDP[8]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_2_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_1_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_0_1_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_0_1_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_1__1_) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_0_1_U6 ( .A1(InverterInxDP[3]), .A2(
        InverterInxDP[5]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_1_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_1_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_0_1_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_0_1_n14), .ZN(
        inverter_gf24_a_mul_b_Xi_mul_Yj_1__0_) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_1_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_0_1_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_0_1_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_0_1_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_1_U3 ( .A(InverterInxDP[3]), .B(
        InverterInxDP[2]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_1_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_1_U2 ( .A(InverterInxDP[5]), .B(
        InverterInxDP[4]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_1_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_0_1_U1 ( .A1(InverterInxDP[2]), .A2(
        InverterInxDP[4]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_1_n13) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_0_U7 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_0_0_n15), .B(
        inverter_gf24_a_mul_b_gf2_mul_0_0_n14), .ZN(
        inverter_gf24_a_mul_b_FFxDN[1]) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_0_0_U6 ( .A1(InverterInxDP[3]), .A2(
        InverterInxDP[1]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_0_n15) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_0_U5 ( .A(
        inverter_gf24_a_mul_b_gf2_mul_0_0_n13), .B(
        inverter_gf24_a_mul_b_gf2_mul_0_0_n14), .ZN(
        inverter_gf24_a_mul_b_FFxDN[0]) );
  NOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_0_U4 ( .A1(
        inverter_gf24_a_mul_b_gf2_mul_0_0_n12), .A2(
        inverter_gf24_a_mul_b_gf2_mul_0_0_n11), .ZN(
        inverter_gf24_a_mul_b_gf2_mul_0_0_n14) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_0_U3 ( .A(InverterInxDP[3]), .B(
        InverterInxDP[2]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_0_n11) );
  XNOR2_X1 inverter_gf24_a_mul_b_gf2_mul_0_0_U2 ( .A(InverterInxDP[1]), .B(
        InverterInxDP[0]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_0_n12) );
  NAND2_X1 inverter_gf24_a_mul_b_gf2_mul_0_0_U1 ( .A1(InverterInxDP[2]), .A2(
        InverterInxDP[0]), .ZN(inverter_gf24_a_mul_b_gf2_mul_0_0_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_U50 ( .A(inverter_gf24_a_mul_e_n64), .B(
        inverter_gf24_a_mul_e_n63), .ZN(InverterOutxD[13]) );
  XNOR2_X1 inverter_gf24_a_mul_e_U49 ( .A(inverter_gf24_a_mul_e_n18), .B(
        inverter_gf24_a_mul_e_n17), .ZN(inverter_gf24_a_mul_e_n63) );
  XOR2_X1 inverter_gf24_a_mul_e_U48 ( .A(inverter_gf24_a_mul_e_n20), .B(
        inverter_gf24_a_mul_e_n19), .Z(inverter_gf24_a_mul_e_n64) );
  XNOR2_X1 inverter_gf24_a_mul_e_U47 ( .A(inverter_gf24_a_mul_e_n62), .B(
        inverter_gf24_a_mul_e_n61), .ZN(InverterOutxD[12]) );
  XNOR2_X1 inverter_gf24_a_mul_e_U46 ( .A(inverter_gf24_a_mul_e_n22), .B(
        inverter_gf24_a_mul_e_n21), .ZN(inverter_gf24_a_mul_e_n61) );
  XOR2_X1 inverter_gf24_a_mul_e_U45 ( .A(inverter_gf24_a_mul_e_n24), .B(
        inverter_gf24_a_mul_e_n23), .Z(inverter_gf24_a_mul_e_n62) );
  XNOR2_X1 inverter_gf24_a_mul_e_U44 ( .A(inverter_gf24_a_mul_e_n60), .B(
        inverter_gf24_a_mul_e_n59), .ZN(InverterOutxD[9]) );
  XNOR2_X1 inverter_gf24_a_mul_e_U43 ( .A(inverter_gf24_a_mul_e_n26), .B(
        inverter_gf24_a_mul_e_n25), .ZN(inverter_gf24_a_mul_e_n59) );
  XOR2_X1 inverter_gf24_a_mul_e_U42 ( .A(inverter_gf24_a_mul_e_n28), .B(
        inverter_gf24_a_mul_e_n27), .Z(inverter_gf24_a_mul_e_n60) );
  XNOR2_X1 inverter_gf24_a_mul_e_U41 ( .A(inverter_gf24_a_mul_e_n58), .B(
        inverter_gf24_a_mul_e_n57), .ZN(InverterOutxD[8]) );
  XNOR2_X1 inverter_gf24_a_mul_e_U40 ( .A(inverter_gf24_a_mul_e_n30), .B(
        inverter_gf24_a_mul_e_n29), .ZN(inverter_gf24_a_mul_e_n57) );
  XOR2_X1 inverter_gf24_a_mul_e_U39 ( .A(inverter_gf24_a_mul_e_n32), .B(
        inverter_gf24_a_mul_e_n31), .Z(inverter_gf24_a_mul_e_n58) );
  XNOR2_X1 inverter_gf24_a_mul_e_U38 ( .A(inverter_gf24_a_mul_e_n56), .B(
        inverter_gf24_a_mul_e_n55), .ZN(InverterOutxD[5]) );
  XNOR2_X1 inverter_gf24_a_mul_e_U37 ( .A(inverter_gf24_a_mul_e_n34), .B(
        inverter_gf24_a_mul_e_n33), .ZN(inverter_gf24_a_mul_e_n55) );
  XOR2_X1 inverter_gf24_a_mul_e_U36 ( .A(inverter_gf24_a_mul_e_n36), .B(
        inverter_gf24_a_mul_e_n35), .Z(inverter_gf24_a_mul_e_n56) );
  XNOR2_X1 inverter_gf24_a_mul_e_U35 ( .A(inverter_gf24_a_mul_e_n54), .B(
        inverter_gf24_a_mul_e_n53), .ZN(InverterOutxD[4]) );
  XNOR2_X1 inverter_gf24_a_mul_e_U34 ( .A(inverter_gf24_a_mul_e_n38), .B(
        inverter_gf24_a_mul_e_n37), .ZN(inverter_gf24_a_mul_e_n53) );
  XOR2_X1 inverter_gf24_a_mul_e_U33 ( .A(inverter_gf24_a_mul_e_n40), .B(
        inverter_gf24_a_mul_e_n39), .Z(inverter_gf24_a_mul_e_n54) );
  XNOR2_X1 inverter_gf24_a_mul_e_U32 ( .A(inverter_gf24_a_mul_e_n52), .B(
        inverter_gf24_a_mul_e_n51), .ZN(InverterOutxD[1]) );
  XNOR2_X1 inverter_gf24_a_mul_e_U31 ( .A(inverter_gf24_a_mul_e_n42), .B(
        inverter_gf24_a_mul_e_n41), .ZN(inverter_gf24_a_mul_e_n51) );
  XOR2_X1 inverter_gf24_a_mul_e_U30 ( .A(inverter_gf24_a_mul_e_n44), .B(
        inverter_gf24_a_mul_e_n43), .Z(inverter_gf24_a_mul_e_n52) );
  XNOR2_X1 inverter_gf24_a_mul_e_U29 ( .A(inverter_gf24_a_mul_e_n50), .B(
        inverter_gf24_a_mul_e_n49), .ZN(InverterOutxD[0]) );
  XNOR2_X1 inverter_gf24_a_mul_e_U28 ( .A(inverter_gf24_a_mul_e_n46), .B(
        inverter_gf24_a_mul_e_n45), .ZN(inverter_gf24_a_mul_e_n49) );
  XOR2_X1 inverter_gf24_a_mul_e_U27 ( .A(inverter_gf24_a_mul_e_n48), .B(
        inverter_gf24_a_mul_e_n47), .Z(inverter_gf24_a_mul_e_n50) );
  XOR2_X1 inverter_gf24_a_mul_e_U26 ( .A(Zinv2xDI[5]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_9__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[19]) );
  XOR2_X1 inverter_gf24_a_mul_e_U25 ( .A(Zinv2xDI[4]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_9__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[18]) );
  XOR2_X1 inverter_gf24_a_mul_e_U24 ( .A(Zinv2xDI[3]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_8__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[17]) );
  XOR2_X1 inverter_gf24_a_mul_e_U23 ( .A(Zinv2xDI[2]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_8__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[16]) );
  XOR2_X1 inverter_gf24_a_mul_e_U22 ( .A(Zinv2xDI[9]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_7__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[15]) );
  XOR2_X1 inverter_gf24_a_mul_e_U21 ( .A(Zinv2xDI[8]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_7__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[14]) );
  XOR2_X1 inverter_gf24_a_mul_e_U20 ( .A(Zinv2xDI[5]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_6__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[13]) );
  XOR2_X1 inverter_gf24_a_mul_e_U19 ( .A(Zinv2xDI[4]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_6__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[12]) );
  XOR2_X1 inverter_gf24_a_mul_e_U18 ( .A(Zinv2xDI[1]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_4__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[9]) );
  XOR2_X1 inverter_gf24_a_mul_e_U17 ( .A(Zinv2xDI[0]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_4__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[8]) );
  XOR2_X1 inverter_gf24_a_mul_e_U16 ( .A(Zinv2xDI[7]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_3__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[7]) );
  XOR2_X1 inverter_gf24_a_mul_e_U15 ( .A(Zinv2xDI[6]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_3__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[6]) );
  XOR2_X1 inverter_gf24_a_mul_e_U14 ( .A(Zinv2xDI[3]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_2__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[5]) );
  XOR2_X1 inverter_gf24_a_mul_e_U13 ( .A(Zinv2xDI[2]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_2__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[4]) );
  XOR2_X1 inverter_gf24_a_mul_e_U12 ( .A(Zinv2xDI[1]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_1__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[3]) );
  XOR2_X1 inverter_gf24_a_mul_e_U11 ( .A(Zinv2xDI[0]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_1__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[2]) );
  XOR2_X1 inverter_gf24_a_mul_e_U10 ( .A(Zinv2xDI[11]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_14__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[29]) );
  XOR2_X1 inverter_gf24_a_mul_e_U9 ( .A(Zinv2xDI[10]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_14__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[28]) );
  XOR2_X1 inverter_gf24_a_mul_e_U8 ( .A(Zinv2xDI[9]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_13__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[27]) );
  XOR2_X1 inverter_gf24_a_mul_e_U7 ( .A(Zinv2xDI[8]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_13__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[26]) );
  XOR2_X1 inverter_gf24_a_mul_e_U6 ( .A(Zinv2xDI[7]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_12__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[25]) );
  XOR2_X1 inverter_gf24_a_mul_e_U5 ( .A(Zinv2xDI[6]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_12__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[24]) );
  XOR2_X1 inverter_gf24_a_mul_e_U4 ( .A(Zinv2xDI[11]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_11__1_), .Z(
        inverter_gf24_a_mul_e_FFxDN[23]) );
  XOR2_X1 inverter_gf24_a_mul_e_U3 ( .A(Zinv2xDI[10]), .B(
        inverter_gf24_a_mul_e_Xi_mul_Yj_11__0_), .Z(
        inverter_gf24_a_mul_e_FFxDN[22]) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_1__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[2]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n48) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_2__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[4]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n45) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_3__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[6]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n46) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_4__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[8]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n39) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_6__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[12]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n37) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_7__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[14]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n38) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_8__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[16]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n29) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_9__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[18]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n30) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_11__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[22]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n32) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_12__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[24]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n23) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_13__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[26]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n24) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_14__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[28]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n21) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_1__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[3]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n44) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_2__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[5]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n41) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_3__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[7]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n42) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_4__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[9]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n35) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_6__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[13]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n33) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_7__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[15]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n34) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_8__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[17]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n25) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_9__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[19]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n26) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_11__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[23]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n28) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_12__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[25]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n19) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_13__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[27]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n20) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_14__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[29]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n17) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_0__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[0]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n47) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_5__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[10]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n40) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_10__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[20]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n31) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_15__0_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[30]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n22) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_0__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[1]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n43) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_5__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[11]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n36) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_10__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[21]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n27) );
  DFF_X1 inverter_gf24_a_mul_e_FFxDP_reg_15__1_ ( .D(
        inverter_gf24_a_mul_e_FFxDN[31]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_a_mul_e_n18) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_3_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_3_3_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_3_3_n14), .ZN(
        inverter_gf24_a_mul_e_FFxDN[31]) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_3_3_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[7]), .A2(inverter_gf24_ExDP_3__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_3_3_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_3_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_3_3_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_3_3_n14), .ZN(
        inverter_gf24_a_mul_e_FFxDN[30]) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_3_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_3_3_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_3_3_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_3_3_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_3_U3 ( .A(
        inverter_gf24_pipelinedAxDP[7]), .B(inverter_gf24_pipelinedAxDP[6]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_3_3_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_3_U2 ( .A(inverter_gf24_ExDP_3__1_), 
        .B(inverter_gf24_ExDP_3__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_3_3_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_3_3_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[6]), .A2(inverter_gf24_ExDP_3__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_3_3_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_2_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_3_2_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_3_2_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_14__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_3_2_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[7]), .A2(inverter_gf24_ExDP_2__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_3_2_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_2_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_3_2_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_3_2_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_14__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_2_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_3_2_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_3_2_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_3_2_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_2_U3 ( .A(
        inverter_gf24_pipelinedAxDP[7]), .B(inverter_gf24_pipelinedAxDP[6]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_3_2_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_2_U2 ( .A(inverter_gf24_ExDP_2__1_), 
        .B(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_3_2_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_3_2_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[6]), .A2(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_3_2_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_1_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_3_1_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_3_1_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_13__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_3_1_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[7]), .A2(inverter_gf24_ExDP_1__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_3_1_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_1_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_3_1_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_3_1_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_13__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_1_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_3_1_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_3_1_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_3_1_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_1_U3 ( .A(
        inverter_gf24_pipelinedAxDP[7]), .B(inverter_gf24_pipelinedAxDP[6]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_3_1_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_1_U2 ( .A(inverter_gf24_ExDP_1__1_), 
        .B(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_3_1_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_3_1_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[6]), .A2(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_3_1_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_0_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_3_0_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_3_0_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_12__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_3_0_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[7]), .A2(inverter_gf24_ExDP_0__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_3_0_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_0_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_3_0_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_3_0_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_12__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_0_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_3_0_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_3_0_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_3_0_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_0_U3 ( .A(
        inverter_gf24_pipelinedAxDP[7]), .B(inverter_gf24_pipelinedAxDP[6]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_3_0_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_3_0_U2 ( .A(inverter_gf24_ExDP_0__1_), 
        .B(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_3_0_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_3_0_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[6]), .A2(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_3_0_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_3_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_2_3_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_2_3_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_11__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_2_3_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[5]), .A2(inverter_gf24_ExDP_3__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_3_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_3_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_2_3_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_2_3_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_11__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_3_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_2_3_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_2_3_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_3_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_3_U3 ( .A(
        inverter_gf24_pipelinedAxDP[5]), .B(inverter_gf24_pipelinedAxDP[4]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_2_3_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_3_U2 ( .A(inverter_gf24_ExDP_3__1_), 
        .B(inverter_gf24_ExDP_3__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_3_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_2_3_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[4]), .A2(inverter_gf24_ExDP_3__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_3_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_2_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n14), .ZN(
        inverter_gf24_a_mul_e_FFxDN[21]) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_2_2_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[5]), .A2(inverter_gf24_ExDP_2__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_2_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n14), .ZN(
        inverter_gf24_a_mul_e_FFxDN[20]) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_2_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_2_U3 ( .A(
        inverter_gf24_pipelinedAxDP[5]), .B(inverter_gf24_pipelinedAxDP[4]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_2_2_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_2_U2 ( .A(inverter_gf24_ExDP_2__1_), 
        .B(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_2_2_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[4]), .A2(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_2_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_1_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_9__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_2_1_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[5]), .A2(inverter_gf24_ExDP_1__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_1_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_9__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_1_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_1_U3 ( .A(
        inverter_gf24_pipelinedAxDP[5]), .B(inverter_gf24_pipelinedAxDP[4]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_2_1_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_1_U2 ( .A(inverter_gf24_ExDP_1__1_), 
        .B(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_2_1_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[4]), .A2(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_1_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_0_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_8__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_2_0_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[5]), .A2(inverter_gf24_ExDP_0__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_0_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_8__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_0_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_0_U3 ( .A(
        inverter_gf24_pipelinedAxDP[5]), .B(inverter_gf24_pipelinedAxDP[4]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_2_0_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_2_0_U2 ( .A(inverter_gf24_ExDP_0__1_), 
        .B(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_2_0_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[4]), .A2(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_2_0_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_3_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_1_3_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_1_3_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_7__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_1_3_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[3]), .A2(inverter_gf24_ExDP_3__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_3_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_3_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_1_3_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_1_3_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_7__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_3_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_1_3_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_1_3_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_3_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_3_U3 ( .A(
        inverter_gf24_pipelinedAxDP[3]), .B(inverter_gf24_pipelinedAxDP[2]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_1_3_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_3_U2 ( .A(inverter_gf24_ExDP_3__1_), 
        .B(inverter_gf24_ExDP_3__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_3_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_1_3_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[2]), .A2(inverter_gf24_ExDP_3__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_3_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_2_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_6__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_1_2_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[3]), .A2(inverter_gf24_ExDP_2__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_2_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_6__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_2_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_2_U3 ( .A(
        inverter_gf24_pipelinedAxDP[3]), .B(inverter_gf24_pipelinedAxDP[2]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_1_2_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_2_U2 ( .A(inverter_gf24_ExDP_2__1_), 
        .B(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_1_2_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[2]), .A2(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_2_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_1_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n14), .ZN(
        inverter_gf24_a_mul_e_FFxDN[11]) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_1_1_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[3]), .A2(inverter_gf24_ExDP_1__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_1_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n14), .ZN(
        inverter_gf24_a_mul_e_FFxDN[10]) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_1_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_1_U3 ( .A(
        inverter_gf24_pipelinedAxDP[3]), .B(inverter_gf24_pipelinedAxDP[2]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_1_1_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_1_U2 ( .A(inverter_gf24_ExDP_1__1_), 
        .B(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_1_1_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[2]), .A2(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_1_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_0_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_4__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_1_0_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[3]), .A2(inverter_gf24_ExDP_0__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_0_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_4__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_0_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_0_U3 ( .A(
        inverter_gf24_pipelinedAxDP[3]), .B(inverter_gf24_pipelinedAxDP[2]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_1_0_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_1_0_U2 ( .A(inverter_gf24_ExDP_0__1_), 
        .B(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_1_0_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[2]), .A2(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_1_0_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_3_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_0_3_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_0_3_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_3__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_0_3_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[1]), .A2(inverter_gf24_ExDP_3__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_3_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_3_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_0_3_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_0_3_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_3__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_3_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_0_3_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_0_3_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_3_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_3_U3 ( .A(
        inverter_gf24_pipelinedAxDP[1]), .B(inverter_gf24_pipelinedAxDP[0]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_0_3_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_3_U2 ( .A(inverter_gf24_ExDP_3__1_), 
        .B(inverter_gf24_ExDP_3__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_3_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_0_3_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[0]), .A2(inverter_gf24_ExDP_3__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_3_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_2_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_2__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_0_2_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[1]), .A2(inverter_gf24_ExDP_2__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_2_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_2__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_2_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_2_U3 ( .A(
        inverter_gf24_pipelinedAxDP[1]), .B(inverter_gf24_pipelinedAxDP[0]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_0_2_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_2_U2 ( .A(inverter_gf24_ExDP_2__1_), 
        .B(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_0_2_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[0]), .A2(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_2_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_1_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_1__1_) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_0_1_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[1]), .A2(inverter_gf24_ExDP_1__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_1_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n14), .ZN(
        inverter_gf24_a_mul_e_Xi_mul_Yj_1__0_) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_1_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_1_U3 ( .A(
        inverter_gf24_pipelinedAxDP[1]), .B(inverter_gf24_pipelinedAxDP[0]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_0_1_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_1_U2 ( .A(inverter_gf24_ExDP_1__1_), 
        .B(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_0_1_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[0]), .A2(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_1_n13) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_0_U7 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n15), .B(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n14), .ZN(
        inverter_gf24_a_mul_e_FFxDN[1]) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_0_0_U6 ( .A1(
        inverter_gf24_pipelinedAxDP[1]), .A2(inverter_gf24_ExDP_0__1_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n15) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_0_U5 ( .A(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n13), .B(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n14), .ZN(
        inverter_gf24_a_mul_e_FFxDN[0]) );
  NOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_0_U4 ( .A1(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n12), .A2(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n11), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n14) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_0_U3 ( .A(
        inverter_gf24_pipelinedAxDP[1]), .B(inverter_gf24_pipelinedAxDP[0]), 
        .ZN(inverter_gf24_a_mul_e_gf2_mul_0_0_n11) );
  XNOR2_X1 inverter_gf24_a_mul_e_gf2_mul_0_0_U2 ( .A(inverter_gf24_ExDP_0__1_), 
        .B(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n12) );
  NAND2_X1 inverter_gf24_a_mul_e_gf2_mul_0_0_U1 ( .A1(
        inverter_gf24_pipelinedAxDP[0]), .A2(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_a_mul_e_gf2_mul_0_0_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_U50 ( .A(inverter_gf24_b_mul_e_n64), .B(
        inverter_gf24_b_mul_e_n63), .ZN(InverterOutxD[15]) );
  XNOR2_X1 inverter_gf24_b_mul_e_U49 ( .A(inverter_gf24_b_mul_e_n18), .B(
        inverter_gf24_b_mul_e_n17), .ZN(inverter_gf24_b_mul_e_n63) );
  XOR2_X1 inverter_gf24_b_mul_e_U48 ( .A(inverter_gf24_b_mul_e_n20), .B(
        inverter_gf24_b_mul_e_n19), .Z(inverter_gf24_b_mul_e_n64) );
  XNOR2_X1 inverter_gf24_b_mul_e_U47 ( .A(inverter_gf24_b_mul_e_n62), .B(
        inverter_gf24_b_mul_e_n61), .ZN(InverterOutxD[14]) );
  XNOR2_X1 inverter_gf24_b_mul_e_U46 ( .A(inverter_gf24_b_mul_e_n22), .B(
        inverter_gf24_b_mul_e_n21), .ZN(inverter_gf24_b_mul_e_n61) );
  XOR2_X1 inverter_gf24_b_mul_e_U45 ( .A(inverter_gf24_b_mul_e_n24), .B(
        inverter_gf24_b_mul_e_n23), .Z(inverter_gf24_b_mul_e_n62) );
  XNOR2_X1 inverter_gf24_b_mul_e_U44 ( .A(inverter_gf24_b_mul_e_n60), .B(
        inverter_gf24_b_mul_e_n59), .ZN(InverterOutxD[11]) );
  XNOR2_X1 inverter_gf24_b_mul_e_U43 ( .A(inverter_gf24_b_mul_e_n26), .B(
        inverter_gf24_b_mul_e_n25), .ZN(inverter_gf24_b_mul_e_n59) );
  XOR2_X1 inverter_gf24_b_mul_e_U42 ( .A(inverter_gf24_b_mul_e_n28), .B(
        inverter_gf24_b_mul_e_n27), .Z(inverter_gf24_b_mul_e_n60) );
  XNOR2_X1 inverter_gf24_b_mul_e_U41 ( .A(inverter_gf24_b_mul_e_n58), .B(
        inverter_gf24_b_mul_e_n57), .ZN(InverterOutxD[10]) );
  XNOR2_X1 inverter_gf24_b_mul_e_U40 ( .A(inverter_gf24_b_mul_e_n30), .B(
        inverter_gf24_b_mul_e_n29), .ZN(inverter_gf24_b_mul_e_n57) );
  XOR2_X1 inverter_gf24_b_mul_e_U39 ( .A(inverter_gf24_b_mul_e_n32), .B(
        inverter_gf24_b_mul_e_n31), .Z(inverter_gf24_b_mul_e_n58) );
  XNOR2_X1 inverter_gf24_b_mul_e_U38 ( .A(inverter_gf24_b_mul_e_n56), .B(
        inverter_gf24_b_mul_e_n55), .ZN(InverterOutxD[7]) );
  XNOR2_X1 inverter_gf24_b_mul_e_U37 ( .A(inverter_gf24_b_mul_e_n34), .B(
        inverter_gf24_b_mul_e_n33), .ZN(inverter_gf24_b_mul_e_n55) );
  XOR2_X1 inverter_gf24_b_mul_e_U36 ( .A(inverter_gf24_b_mul_e_n36), .B(
        inverter_gf24_b_mul_e_n35), .Z(inverter_gf24_b_mul_e_n56) );
  XNOR2_X1 inverter_gf24_b_mul_e_U35 ( .A(inverter_gf24_b_mul_e_n54), .B(
        inverter_gf24_b_mul_e_n53), .ZN(InverterOutxD[6]) );
  XNOR2_X1 inverter_gf24_b_mul_e_U34 ( .A(inverter_gf24_b_mul_e_n38), .B(
        inverter_gf24_b_mul_e_n37), .ZN(inverter_gf24_b_mul_e_n53) );
  XOR2_X1 inverter_gf24_b_mul_e_U33 ( .A(inverter_gf24_b_mul_e_n40), .B(
        inverter_gf24_b_mul_e_n39), .Z(inverter_gf24_b_mul_e_n54) );
  XNOR2_X1 inverter_gf24_b_mul_e_U32 ( .A(inverter_gf24_b_mul_e_n52), .B(
        inverter_gf24_b_mul_e_n51), .ZN(InverterOutxD[3]) );
  XNOR2_X1 inverter_gf24_b_mul_e_U31 ( .A(inverter_gf24_b_mul_e_n42), .B(
        inverter_gf24_b_mul_e_n41), .ZN(inverter_gf24_b_mul_e_n51) );
  XOR2_X1 inverter_gf24_b_mul_e_U30 ( .A(inverter_gf24_b_mul_e_n44), .B(
        inverter_gf24_b_mul_e_n43), .Z(inverter_gf24_b_mul_e_n52) );
  XNOR2_X1 inverter_gf24_b_mul_e_U29 ( .A(inverter_gf24_b_mul_e_n50), .B(
        inverter_gf24_b_mul_e_n49), .ZN(InverterOutxD[2]) );
  XNOR2_X1 inverter_gf24_b_mul_e_U28 ( .A(inverter_gf24_b_mul_e_n46), .B(
        inverter_gf24_b_mul_e_n45), .ZN(inverter_gf24_b_mul_e_n49) );
  XOR2_X1 inverter_gf24_b_mul_e_U27 ( .A(inverter_gf24_b_mul_e_n48), .B(
        inverter_gf24_b_mul_e_n47), .Z(inverter_gf24_b_mul_e_n50) );
  XOR2_X1 inverter_gf24_b_mul_e_U26 ( .A(Zinv3xDI[5]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_9__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[19]) );
  XOR2_X1 inverter_gf24_b_mul_e_U25 ( .A(Zinv3xDI[4]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_9__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[18]) );
  XOR2_X1 inverter_gf24_b_mul_e_U24 ( .A(Zinv3xDI[3]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_8__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[17]) );
  XOR2_X1 inverter_gf24_b_mul_e_U23 ( .A(Zinv3xDI[2]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_8__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[16]) );
  XOR2_X1 inverter_gf24_b_mul_e_U22 ( .A(Zinv3xDI[9]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_7__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[15]) );
  XOR2_X1 inverter_gf24_b_mul_e_U21 ( .A(Zinv3xDI[8]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_7__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[14]) );
  XOR2_X1 inverter_gf24_b_mul_e_U20 ( .A(Zinv3xDI[5]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_6__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[13]) );
  XOR2_X1 inverter_gf24_b_mul_e_U19 ( .A(Zinv3xDI[4]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_6__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[12]) );
  XOR2_X1 inverter_gf24_b_mul_e_U18 ( .A(Zinv3xDI[1]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_4__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[9]) );
  XOR2_X1 inverter_gf24_b_mul_e_U17 ( .A(Zinv3xDI[0]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_4__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[8]) );
  XOR2_X1 inverter_gf24_b_mul_e_U16 ( .A(Zinv3xDI[7]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_3__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[7]) );
  XOR2_X1 inverter_gf24_b_mul_e_U15 ( .A(Zinv3xDI[6]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_3__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[6]) );
  XOR2_X1 inverter_gf24_b_mul_e_U14 ( .A(Zinv3xDI[3]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_2__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[5]) );
  XOR2_X1 inverter_gf24_b_mul_e_U13 ( .A(Zinv3xDI[2]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_2__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[4]) );
  XOR2_X1 inverter_gf24_b_mul_e_U12 ( .A(Zinv3xDI[1]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_1__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[3]) );
  XOR2_X1 inverter_gf24_b_mul_e_U11 ( .A(Zinv3xDI[0]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_1__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[2]) );
  XOR2_X1 inverter_gf24_b_mul_e_U10 ( .A(Zinv3xDI[11]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_14__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[29]) );
  XOR2_X1 inverter_gf24_b_mul_e_U9 ( .A(Zinv3xDI[10]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_14__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[28]) );
  XOR2_X1 inverter_gf24_b_mul_e_U8 ( .A(Zinv3xDI[9]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_13__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[27]) );
  XOR2_X1 inverter_gf24_b_mul_e_U7 ( .A(Zinv3xDI[8]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_13__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[26]) );
  XOR2_X1 inverter_gf24_b_mul_e_U6 ( .A(Zinv3xDI[7]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_12__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[25]) );
  XOR2_X1 inverter_gf24_b_mul_e_U5 ( .A(Zinv3xDI[6]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_12__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[24]) );
  XOR2_X1 inverter_gf24_b_mul_e_U4 ( .A(Zinv3xDI[11]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_11__1_), .Z(
        inverter_gf24_b_mul_e_FFxDN[23]) );
  XOR2_X1 inverter_gf24_b_mul_e_U3 ( .A(Zinv3xDI[10]), .B(
        inverter_gf24_b_mul_e_Xi_mul_Yj_11__0_), .Z(
        inverter_gf24_b_mul_e_FFxDN[22]) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_1__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[2]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n48) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_2__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[4]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n45) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_3__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[6]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n46) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_4__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[8]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n39) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_6__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[12]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n37) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_7__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[14]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n38) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_8__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[16]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n29) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_9__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[18]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n30) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_11__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[22]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n32) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_12__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[24]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n23) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_13__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[26]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n24) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_14__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[28]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n21) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_1__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[3]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n44) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_2__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[5]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n41) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_3__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[7]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n42) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_4__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[9]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n35) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_6__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[13]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n33) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_7__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[15]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n34) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_8__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[17]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n25) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_9__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[19]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n26) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_11__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[23]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n28) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_12__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[25]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n19) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_13__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[27]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n20) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_14__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[29]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n17) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_0__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[0]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n47) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_5__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[10]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n40) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_10__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[20]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n31) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_15__0_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[30]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n22) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_0__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[1]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n43) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_5__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[11]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n36) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_10__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[21]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n27) );
  DFF_X1 inverter_gf24_b_mul_e_FFxDP_reg_15__1_ ( .D(
        inverter_gf24_b_mul_e_FFxDN[31]), .CK(ClkxCI), .Q(), .QN(
        inverter_gf24_b_mul_e_n18) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_3_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_3_3_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_3_3_n14), .ZN(
        inverter_gf24_b_mul_e_FFxDN[31]) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_3_3_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[7]), .A2(inverter_gf24_ExDP_3__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_3_3_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_3_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_3_3_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_3_3_n14), .ZN(
        inverter_gf24_b_mul_e_FFxDN[30]) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_3_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_3_3_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_3_3_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_3_3_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_3_U3 ( .A(
        inverter_gf24_pipelinedBxDP[7]), .B(inverter_gf24_pipelinedBxDP[6]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_3_3_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_3_U2 ( .A(inverter_gf24_ExDP_3__1_), 
        .B(inverter_gf24_ExDP_3__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_3_3_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_3_3_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[6]), .A2(inverter_gf24_ExDP_3__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_3_3_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_2_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_3_2_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_3_2_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_14__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_3_2_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[7]), .A2(inverter_gf24_ExDP_2__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_3_2_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_2_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_3_2_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_3_2_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_14__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_2_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_3_2_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_3_2_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_3_2_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_2_U3 ( .A(
        inverter_gf24_pipelinedBxDP[7]), .B(inverter_gf24_pipelinedBxDP[6]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_3_2_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_2_U2 ( .A(inverter_gf24_ExDP_2__1_), 
        .B(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_3_2_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_3_2_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[6]), .A2(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_3_2_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_1_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_3_1_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_3_1_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_13__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_3_1_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[7]), .A2(inverter_gf24_ExDP_1__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_3_1_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_1_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_3_1_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_3_1_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_13__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_1_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_3_1_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_3_1_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_3_1_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_1_U3 ( .A(
        inverter_gf24_pipelinedBxDP[7]), .B(inverter_gf24_pipelinedBxDP[6]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_3_1_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_1_U2 ( .A(inverter_gf24_ExDP_1__1_), 
        .B(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_3_1_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_3_1_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[6]), .A2(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_3_1_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_0_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_3_0_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_3_0_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_12__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_3_0_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[7]), .A2(inverter_gf24_ExDP_0__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_3_0_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_0_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_3_0_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_3_0_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_12__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_0_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_3_0_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_3_0_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_3_0_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_0_U3 ( .A(
        inverter_gf24_pipelinedBxDP[7]), .B(inverter_gf24_pipelinedBxDP[6]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_3_0_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_3_0_U2 ( .A(inverter_gf24_ExDP_0__1_), 
        .B(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_3_0_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_3_0_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[6]), .A2(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_3_0_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_3_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_2_3_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_2_3_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_11__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_2_3_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[5]), .A2(inverter_gf24_ExDP_3__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_3_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_3_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_2_3_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_2_3_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_11__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_3_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_2_3_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_2_3_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_3_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_3_U3 ( .A(
        inverter_gf24_pipelinedBxDP[5]), .B(inverter_gf24_pipelinedBxDP[4]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_2_3_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_3_U2 ( .A(inverter_gf24_ExDP_3__1_), 
        .B(inverter_gf24_ExDP_3__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_3_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_2_3_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[4]), .A2(inverter_gf24_ExDP_3__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_3_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_2_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n14), .ZN(
        inverter_gf24_b_mul_e_FFxDN[21]) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_2_2_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[5]), .A2(inverter_gf24_ExDP_2__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_2_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n14), .ZN(
        inverter_gf24_b_mul_e_FFxDN[20]) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_2_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_2_U3 ( .A(
        inverter_gf24_pipelinedBxDP[5]), .B(inverter_gf24_pipelinedBxDP[4]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_2_2_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_2_U2 ( .A(inverter_gf24_ExDP_2__1_), 
        .B(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_2_2_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[4]), .A2(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_2_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_1_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_9__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_2_1_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[5]), .A2(inverter_gf24_ExDP_1__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_1_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_9__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_1_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_1_U3 ( .A(
        inverter_gf24_pipelinedBxDP[5]), .B(inverter_gf24_pipelinedBxDP[4]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_2_1_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_1_U2 ( .A(inverter_gf24_ExDP_1__1_), 
        .B(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_2_1_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[4]), .A2(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_1_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_0_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_8__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_2_0_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[5]), .A2(inverter_gf24_ExDP_0__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_0_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_8__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_0_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_0_U3 ( .A(
        inverter_gf24_pipelinedBxDP[5]), .B(inverter_gf24_pipelinedBxDP[4]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_2_0_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_2_0_U2 ( .A(inverter_gf24_ExDP_0__1_), 
        .B(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_2_0_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[4]), .A2(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_2_0_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_3_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_1_3_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_1_3_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_7__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_1_3_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[3]), .A2(inverter_gf24_ExDP_3__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_3_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_3_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_1_3_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_1_3_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_7__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_3_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_1_3_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_1_3_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_3_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_3_U3 ( .A(
        inverter_gf24_pipelinedBxDP[3]), .B(inverter_gf24_pipelinedBxDP[2]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_1_3_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_3_U2 ( .A(inverter_gf24_ExDP_3__1_), 
        .B(inverter_gf24_ExDP_3__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_3_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_1_3_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[2]), .A2(inverter_gf24_ExDP_3__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_3_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_2_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_6__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_1_2_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[3]), .A2(inverter_gf24_ExDP_2__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_2_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_6__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_2_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_2_U3 ( .A(
        inverter_gf24_pipelinedBxDP[3]), .B(inverter_gf24_pipelinedBxDP[2]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_1_2_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_2_U2 ( .A(inverter_gf24_ExDP_2__1_), 
        .B(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_1_2_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[2]), .A2(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_2_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_1_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n14), .ZN(
        inverter_gf24_b_mul_e_FFxDN[11]) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_1_1_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[3]), .A2(inverter_gf24_ExDP_1__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_1_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n14), .ZN(
        inverter_gf24_b_mul_e_FFxDN[10]) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_1_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_1_U3 ( .A(
        inverter_gf24_pipelinedBxDP[3]), .B(inverter_gf24_pipelinedBxDP[2]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_1_1_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_1_U2 ( .A(inverter_gf24_ExDP_1__1_), 
        .B(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_1_1_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[2]), .A2(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_1_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_0_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_4__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_1_0_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[3]), .A2(inverter_gf24_ExDP_0__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_0_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_4__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_0_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_0_U3 ( .A(
        inverter_gf24_pipelinedBxDP[3]), .B(inverter_gf24_pipelinedBxDP[2]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_1_0_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_1_0_U2 ( .A(inverter_gf24_ExDP_0__1_), 
        .B(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_1_0_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[2]), .A2(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_1_0_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_3_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_0_3_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_0_3_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_3__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_0_3_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[1]), .A2(inverter_gf24_ExDP_3__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_3_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_3_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_0_3_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_0_3_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_3__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_3_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_0_3_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_0_3_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_3_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_3_U3 ( .A(
        inverter_gf24_pipelinedBxDP[1]), .B(inverter_gf24_pipelinedBxDP[0]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_0_3_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_3_U2 ( .A(inverter_gf24_ExDP_3__1_), 
        .B(inverter_gf24_ExDP_3__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_3_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_0_3_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[0]), .A2(inverter_gf24_ExDP_3__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_3_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_2_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_2__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_0_2_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[1]), .A2(inverter_gf24_ExDP_2__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_2_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_2__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_2_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_2_U3 ( .A(
        inverter_gf24_pipelinedBxDP[1]), .B(inverter_gf24_pipelinedBxDP[0]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_0_2_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_2_U2 ( .A(inverter_gf24_ExDP_2__1_), 
        .B(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_0_2_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[0]), .A2(inverter_gf24_ExDP_2__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_2_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_1_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_1__1_) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_0_1_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[1]), .A2(inverter_gf24_ExDP_1__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_1_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n14), .ZN(
        inverter_gf24_b_mul_e_Xi_mul_Yj_1__0_) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_1_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_1_U3 ( .A(
        inverter_gf24_pipelinedBxDP[1]), .B(inverter_gf24_pipelinedBxDP[0]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_0_1_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_1_U2 ( .A(inverter_gf24_ExDP_1__1_), 
        .B(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_0_1_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[0]), .A2(inverter_gf24_ExDP_1__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_1_n13) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_0_U7 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n15), .B(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n14), .ZN(
        inverter_gf24_b_mul_e_FFxDN[1]) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_0_0_U6 ( .A1(
        inverter_gf24_pipelinedBxDP[1]), .A2(inverter_gf24_ExDP_0__1_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n15) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_0_U5 ( .A(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n13), .B(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n14), .ZN(
        inverter_gf24_b_mul_e_FFxDN[0]) );
  NOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_0_U4 ( .A1(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n12), .A2(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n11), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n14) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_0_U3 ( .A(
        inverter_gf24_pipelinedBxDP[1]), .B(inverter_gf24_pipelinedBxDP[0]), 
        .ZN(inverter_gf24_b_mul_e_gf2_mul_0_0_n11) );
  XNOR2_X1 inverter_gf24_b_mul_e_gf2_mul_0_0_U2 ( .A(inverter_gf24_ExDP_0__1_), 
        .B(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n12) );
  NAND2_X1 inverter_gf24_b_mul_e_gf2_mul_0_0_U1 ( .A1(
        inverter_gf24_pipelinedBxDP[0]), .A2(inverter_gf24_ExDP_0__0_), .ZN(
        inverter_gf24_b_mul_e_gf2_mul_0_0_n13) );
  XNOR2_X1 mult_msb_U98 ( .A(mult_msb_n128), .B(mult_msb_n127), .ZN(
        InvUnmappedxD[31]) );
  XNOR2_X1 mult_msb_U97 ( .A(mult_msb_n34), .B(mult_msb_n33), .ZN(
        mult_msb_n127) );
  XOR2_X1 mult_msb_U96 ( .A(mult_msb_n36), .B(mult_msb_n35), .Z(mult_msb_n128)
         );
  XNOR2_X1 mult_msb_U95 ( .A(mult_msb_n126), .B(mult_msb_n125), .ZN(
        InvUnmappedxD[30]) );
  XNOR2_X1 mult_msb_U94 ( .A(mult_msb_n38), .B(mult_msb_n37), .ZN(
        mult_msb_n125) );
  XOR2_X1 mult_msb_U93 ( .A(mult_msb_n40), .B(mult_msb_n39), .Z(mult_msb_n126)
         );
  XNOR2_X1 mult_msb_U92 ( .A(mult_msb_n124), .B(mult_msb_n123), .ZN(
        InvUnmappedxD[29]) );
  XNOR2_X1 mult_msb_U91 ( .A(mult_msb_n42), .B(mult_msb_n41), .ZN(
        mult_msb_n123) );
  XOR2_X1 mult_msb_U90 ( .A(mult_msb_n44), .B(mult_msb_n43), .Z(mult_msb_n124)
         );
  XNOR2_X1 mult_msb_U89 ( .A(mult_msb_n122), .B(mult_msb_n121), .ZN(
        InvUnmappedxD[28]) );
  XNOR2_X1 mult_msb_U88 ( .A(mult_msb_n46), .B(mult_msb_n45), .ZN(
        mult_msb_n121) );
  XOR2_X1 mult_msb_U87 ( .A(mult_msb_n48), .B(mult_msb_n47), .Z(mult_msb_n122)
         );
  XNOR2_X1 mult_msb_U86 ( .A(mult_msb_n120), .B(mult_msb_n119), .ZN(
        InvUnmappedxD[23]) );
  XNOR2_X1 mult_msb_U85 ( .A(mult_msb_n50), .B(mult_msb_n49), .ZN(
        mult_msb_n119) );
  XOR2_X1 mult_msb_U84 ( .A(mult_msb_n52), .B(mult_msb_n51), .Z(mult_msb_n120)
         );
  XNOR2_X1 mult_msb_U83 ( .A(mult_msb_n118), .B(mult_msb_n117), .ZN(
        InvUnmappedxD[22]) );
  XNOR2_X1 mult_msb_U82 ( .A(mult_msb_n54), .B(mult_msb_n53), .ZN(
        mult_msb_n117) );
  XOR2_X1 mult_msb_U81 ( .A(mult_msb_n56), .B(mult_msb_n55), .Z(mult_msb_n118)
         );
  XNOR2_X1 mult_msb_U80 ( .A(mult_msb_n116), .B(mult_msb_n115), .ZN(
        InvUnmappedxD[21]) );
  XNOR2_X1 mult_msb_U79 ( .A(mult_msb_n58), .B(mult_msb_n57), .ZN(
        mult_msb_n115) );
  XOR2_X1 mult_msb_U78 ( .A(mult_msb_n60), .B(mult_msb_n59), .Z(mult_msb_n116)
         );
  XNOR2_X1 mult_msb_U77 ( .A(mult_msb_n114), .B(mult_msb_n113), .ZN(
        InvUnmappedxD[20]) );
  XNOR2_X1 mult_msb_U76 ( .A(mult_msb_n62), .B(mult_msb_n61), .ZN(
        mult_msb_n113) );
  XOR2_X1 mult_msb_U75 ( .A(mult_msb_n64), .B(mult_msb_n63), .Z(mult_msb_n114)
         );
  XNOR2_X1 mult_msb_U74 ( .A(mult_msb_n112), .B(mult_msb_n111), .ZN(
        InvUnmappedxD[15]) );
  XNOR2_X1 mult_msb_U73 ( .A(mult_msb_n66), .B(mult_msb_n65), .ZN(
        mult_msb_n111) );
  XOR2_X1 mult_msb_U72 ( .A(mult_msb_n68), .B(mult_msb_n67), .Z(mult_msb_n112)
         );
  XNOR2_X1 mult_msb_U71 ( .A(mult_msb_n110), .B(mult_msb_n109), .ZN(
        InvUnmappedxD[14]) );
  XNOR2_X1 mult_msb_U70 ( .A(mult_msb_n70), .B(mult_msb_n69), .ZN(
        mult_msb_n109) );
  XOR2_X1 mult_msb_U69 ( .A(mult_msb_n72), .B(mult_msb_n71), .Z(mult_msb_n110)
         );
  XNOR2_X1 mult_msb_U68 ( .A(mult_msb_n108), .B(mult_msb_n107), .ZN(
        InvUnmappedxD[13]) );
  XNOR2_X1 mult_msb_U67 ( .A(mult_msb_n74), .B(mult_msb_n73), .ZN(
        mult_msb_n107) );
  XOR2_X1 mult_msb_U66 ( .A(mult_msb_n76), .B(mult_msb_n75), .Z(mult_msb_n108)
         );
  XNOR2_X1 mult_msb_U65 ( .A(mult_msb_n106), .B(mult_msb_n105), .ZN(
        InvUnmappedxD[12]) );
  XNOR2_X1 mult_msb_U64 ( .A(mult_msb_n78), .B(mult_msb_n77), .ZN(
        mult_msb_n105) );
  XOR2_X1 mult_msb_U63 ( .A(mult_msb_n80), .B(mult_msb_n79), .Z(mult_msb_n106)
         );
  XNOR2_X1 mult_msb_U62 ( .A(mult_msb_n104), .B(mult_msb_n103), .ZN(
        InvUnmappedxD[7]) );
  XNOR2_X1 mult_msb_U61 ( .A(mult_msb_n82), .B(mult_msb_n81), .ZN(
        mult_msb_n103) );
  XOR2_X1 mult_msb_U60 ( .A(mult_msb_n84), .B(mult_msb_n83), .Z(mult_msb_n104)
         );
  XNOR2_X1 mult_msb_U59 ( .A(mult_msb_n102), .B(mult_msb_n101), .ZN(
        InvUnmappedxD[6]) );
  XNOR2_X1 mult_msb_U58 ( .A(mult_msb_n86), .B(mult_msb_n85), .ZN(
        mult_msb_n101) );
  XOR2_X1 mult_msb_U57 ( .A(mult_msb_n88), .B(mult_msb_n87), .Z(mult_msb_n102)
         );
  XNOR2_X1 mult_msb_U56 ( .A(mult_msb_n100), .B(mult_msb_n99), .ZN(
        InvUnmappedxD[5]) );
  XNOR2_X1 mult_msb_U55 ( .A(mult_msb_n90), .B(mult_msb_n89), .ZN(mult_msb_n99) );
  XOR2_X1 mult_msb_U54 ( .A(mult_msb_n92), .B(mult_msb_n91), .Z(mult_msb_n100)
         );
  XNOR2_X1 mult_msb_U53 ( .A(mult_msb_n98), .B(mult_msb_n97), .ZN(
        InvUnmappedxD[4]) );
  XNOR2_X1 mult_msb_U52 ( .A(mult_msb_n94), .B(mult_msb_n93), .ZN(mult_msb_n97) );
  XOR2_X1 mult_msb_U51 ( .A(mult_msb_n96), .B(mult_msb_n95), .Z(mult_msb_n98)
         );
  XOR2_X1 mult_msb_U50 ( .A(Zmul2xDI[11]), .B(mult_msb_Xi_mul_Yj_9__3_), .Z(
        mult_msb_FFxDN[39]) );
  XOR2_X1 mult_msb_U49 ( .A(Zmul2xDI[10]), .B(mult_msb_Xi_mul_Yj_9__2_), .Z(
        mult_msb_FFxDN[38]) );
  XOR2_X1 mult_msb_U48 ( .A(Zmul2xDI[9]), .B(mult_msb_Xi_mul_Yj_9__1_), .Z(
        mult_msb_FFxDN[37]) );
  XOR2_X1 mult_msb_U47 ( .A(Zmul2xDI[8]), .B(mult_msb_Xi_mul_Yj_9__0_), .Z(
        mult_msb_FFxDN[36]) );
  XOR2_X1 mult_msb_U46 ( .A(Zmul2xDI[7]), .B(mult_msb_Xi_mul_Yj_8__3_), .Z(
        mult_msb_FFxDN[35]) );
  XOR2_X1 mult_msb_U45 ( .A(Zmul2xDI[6]), .B(mult_msb_Xi_mul_Yj_8__2_), .Z(
        mult_msb_FFxDN[34]) );
  XOR2_X1 mult_msb_U44 ( .A(Zmul2xDI[5]), .B(mult_msb_Xi_mul_Yj_8__1_), .Z(
        mult_msb_FFxDN[33]) );
  XOR2_X1 mult_msb_U43 ( .A(Zmul2xDI[4]), .B(mult_msb_Xi_mul_Yj_8__0_), .Z(
        mult_msb_FFxDN[32]) );
  XOR2_X1 mult_msb_U42 ( .A(Zmul2xDI[19]), .B(mult_msb_Xi_mul_Yj_7__3_), .Z(
        mult_msb_FFxDN[31]) );
  XOR2_X1 mult_msb_U41 ( .A(Zmul2xDI[18]), .B(mult_msb_Xi_mul_Yj_7__2_), .Z(
        mult_msb_FFxDN[30]) );
  XOR2_X1 mult_msb_U40 ( .A(Zmul2xDI[17]), .B(mult_msb_Xi_mul_Yj_7__1_), .Z(
        mult_msb_FFxDN[29]) );
  XOR2_X1 mult_msb_U39 ( .A(Zmul2xDI[16]), .B(mult_msb_Xi_mul_Yj_7__0_), .Z(
        mult_msb_FFxDN[28]) );
  XOR2_X1 mult_msb_U38 ( .A(Zmul2xDI[11]), .B(mult_msb_Xi_mul_Yj_6__3_), .Z(
        mult_msb_FFxDN[27]) );
  XOR2_X1 mult_msb_U37 ( .A(Zmul2xDI[10]), .B(mult_msb_Xi_mul_Yj_6__2_), .Z(
        mult_msb_FFxDN[26]) );
  XOR2_X1 mult_msb_U36 ( .A(Zmul2xDI[9]), .B(mult_msb_Xi_mul_Yj_6__1_), .Z(
        mult_msb_FFxDN[25]) );
  XOR2_X1 mult_msb_U35 ( .A(Zmul2xDI[8]), .B(mult_msb_Xi_mul_Yj_6__0_), .Z(
        mult_msb_FFxDN[24]) );
  XOR2_X1 mult_msb_U34 ( .A(Zmul2xDI[3]), .B(mult_msb_Xi_mul_Yj_4__3_), .Z(
        mult_msb_FFxDN[19]) );
  XOR2_X1 mult_msb_U33 ( .A(Zmul2xDI[2]), .B(mult_msb_Xi_mul_Yj_4__2_), .Z(
        mult_msb_FFxDN[18]) );
  XOR2_X1 mult_msb_U32 ( .A(Zmul2xDI[1]), .B(mult_msb_Xi_mul_Yj_4__1_), .Z(
        mult_msb_FFxDN[17]) );
  XOR2_X1 mult_msb_U31 ( .A(Zmul2xDI[0]), .B(mult_msb_Xi_mul_Yj_4__0_), .Z(
        mult_msb_FFxDN[16]) );
  XOR2_X1 mult_msb_U30 ( .A(Zmul2xDI[15]), .B(mult_msb_Xi_mul_Yj_3__3_), .Z(
        mult_msb_FFxDN[15]) );
  XOR2_X1 mult_msb_U29 ( .A(Zmul2xDI[14]), .B(mult_msb_Xi_mul_Yj_3__2_), .Z(
        mult_msb_FFxDN[14]) );
  XOR2_X1 mult_msb_U28 ( .A(Zmul2xDI[13]), .B(mult_msb_Xi_mul_Yj_3__1_), .Z(
        mult_msb_FFxDN[13]) );
  XOR2_X1 mult_msb_U27 ( .A(Zmul2xDI[12]), .B(mult_msb_Xi_mul_Yj_3__0_), .Z(
        mult_msb_FFxDN[12]) );
  XOR2_X1 mult_msb_U26 ( .A(Zmul2xDI[7]), .B(mult_msb_Xi_mul_Yj_2__3_), .Z(
        mult_msb_FFxDN[11]) );
  XOR2_X1 mult_msb_U25 ( .A(Zmul2xDI[6]), .B(mult_msb_Xi_mul_Yj_2__2_), .Z(
        mult_msb_FFxDN[10]) );
  XOR2_X1 mult_msb_U24 ( .A(Zmul2xDI[5]), .B(mult_msb_Xi_mul_Yj_2__1_), .Z(
        mult_msb_FFxDN[9]) );
  XOR2_X1 mult_msb_U23 ( .A(Zmul2xDI[4]), .B(mult_msb_Xi_mul_Yj_2__0_), .Z(
        mult_msb_FFxDN[8]) );
  XOR2_X1 mult_msb_U22 ( .A(Zmul2xDI[3]), .B(mult_msb_Xi_mul_Yj_1__3_), .Z(
        mult_msb_FFxDN[7]) );
  XOR2_X1 mult_msb_U21 ( .A(Zmul2xDI[2]), .B(mult_msb_Xi_mul_Yj_1__2_), .Z(
        mult_msb_FFxDN[6]) );
  XOR2_X1 mult_msb_U20 ( .A(Zmul2xDI[1]), .B(mult_msb_Xi_mul_Yj_1__1_), .Z(
        mult_msb_FFxDN[5]) );
  XOR2_X1 mult_msb_U19 ( .A(Zmul2xDI[0]), .B(mult_msb_Xi_mul_Yj_1__0_), .Z(
        mult_msb_FFxDN[4]) );
  XOR2_X1 mult_msb_U18 ( .A(Zmul2xDI[23]), .B(mult_msb_Xi_mul_Yj_14__3_), .Z(
        mult_msb_FFxDN[59]) );
  XOR2_X1 mult_msb_U17 ( .A(Zmul2xDI[22]), .B(mult_msb_Xi_mul_Yj_14__2_), .Z(
        mult_msb_FFxDN[58]) );
  XOR2_X1 mult_msb_U16 ( .A(Zmul2xDI[21]), .B(mult_msb_Xi_mul_Yj_14__1_), .Z(
        mult_msb_FFxDN[57]) );
  XOR2_X1 mult_msb_U15 ( .A(Zmul2xDI[20]), .B(mult_msb_Xi_mul_Yj_14__0_), .Z(
        mult_msb_FFxDN[56]) );
  XOR2_X1 mult_msb_U14 ( .A(Zmul2xDI[19]), .B(mult_msb_Xi_mul_Yj_13__3_), .Z(
        mult_msb_FFxDN[55]) );
  XOR2_X1 mult_msb_U13 ( .A(Zmul2xDI[18]), .B(mult_msb_Xi_mul_Yj_13__2_), .Z(
        mult_msb_FFxDN[54]) );
  XOR2_X1 mult_msb_U12 ( .A(Zmul2xDI[17]), .B(mult_msb_Xi_mul_Yj_13__1_), .Z(
        mult_msb_FFxDN[53]) );
  XOR2_X1 mult_msb_U11 ( .A(Zmul2xDI[16]), .B(mult_msb_Xi_mul_Yj_13__0_), .Z(
        mult_msb_FFxDN[52]) );
  XOR2_X1 mult_msb_U10 ( .A(Zmul2xDI[15]), .B(mult_msb_Xi_mul_Yj_12__3_), .Z(
        mult_msb_FFxDN[51]) );
  XOR2_X1 mult_msb_U9 ( .A(Zmul2xDI[14]), .B(mult_msb_Xi_mul_Yj_12__2_), .Z(
        mult_msb_FFxDN[50]) );
  XOR2_X1 mult_msb_U8 ( .A(Zmul2xDI[13]), .B(mult_msb_Xi_mul_Yj_12__1_), .Z(
        mult_msb_FFxDN[49]) );
  XOR2_X1 mult_msb_U7 ( .A(Zmul2xDI[12]), .B(mult_msb_Xi_mul_Yj_12__0_), .Z(
        mult_msb_FFxDN[48]) );
  XOR2_X1 mult_msb_U6 ( .A(Zmul2xDI[23]), .B(mult_msb_Xi_mul_Yj_11__3_), .Z(
        mult_msb_FFxDN[47]) );
  XOR2_X1 mult_msb_U5 ( .A(Zmul2xDI[22]), .B(mult_msb_Xi_mul_Yj_11__2_), .Z(
        mult_msb_FFxDN[46]) );
  XOR2_X1 mult_msb_U4 ( .A(Zmul2xDI[21]), .B(mult_msb_Xi_mul_Yj_11__1_), .Z(
        mult_msb_FFxDN[45]) );
  XOR2_X1 mult_msb_U3 ( .A(Zmul2xDI[20]), .B(mult_msb_Xi_mul_Yj_11__0_), .Z(
        mult_msb_FFxDN[44]) );
  DFF_X1 mult_msb_FFxDP_reg_1__3_ ( .D(mult_msb_FFxDN[7]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n84) );
  DFF_X1 mult_msb_FFxDP_reg_2__3_ ( .D(mult_msb_FFxDN[11]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n81) );
  DFF_X1 mult_msb_FFxDP_reg_3__3_ ( .D(mult_msb_FFxDN[15]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n82) );
  DFF_X1 mult_msb_FFxDP_reg_4__3_ ( .D(mult_msb_FFxDN[19]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n67) );
  DFF_X1 mult_msb_FFxDP_reg_6__3_ ( .D(mult_msb_FFxDN[27]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n65) );
  DFF_X1 mult_msb_FFxDP_reg_7__3_ ( .D(mult_msb_FFxDN[31]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n66) );
  DFF_X1 mult_msb_FFxDP_reg_8__3_ ( .D(mult_msb_FFxDN[35]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n49) );
  DFF_X1 mult_msb_FFxDP_reg_9__3_ ( .D(mult_msb_FFxDN[39]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n50) );
  DFF_X1 mult_msb_FFxDP_reg_11__3_ ( .D(mult_msb_FFxDN[47]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n52) );
  DFF_X1 mult_msb_FFxDP_reg_12__3_ ( .D(mult_msb_FFxDN[51]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n35) );
  DFF_X1 mult_msb_FFxDP_reg_13__3_ ( .D(mult_msb_FFxDN[55]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n36) );
  DFF_X1 mult_msb_FFxDP_reg_14__3_ ( .D(mult_msb_FFxDN[59]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n33) );
  DFF_X1 mult_msb_FFxDP_reg_1__1_ ( .D(mult_msb_FFxDN[5]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n92) );
  DFF_X1 mult_msb_FFxDP_reg_2__1_ ( .D(mult_msb_FFxDN[9]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n89) );
  DFF_X1 mult_msb_FFxDP_reg_3__1_ ( .D(mult_msb_FFxDN[13]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n90) );
  DFF_X1 mult_msb_FFxDP_reg_4__1_ ( .D(mult_msb_FFxDN[17]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n75) );
  DFF_X1 mult_msb_FFxDP_reg_6__1_ ( .D(mult_msb_FFxDN[25]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n73) );
  DFF_X1 mult_msb_FFxDP_reg_7__1_ ( .D(mult_msb_FFxDN[29]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n74) );
  DFF_X1 mult_msb_FFxDP_reg_8__1_ ( .D(mult_msb_FFxDN[33]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n57) );
  DFF_X1 mult_msb_FFxDP_reg_9__1_ ( .D(mult_msb_FFxDN[37]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n58) );
  DFF_X1 mult_msb_FFxDP_reg_11__1_ ( .D(mult_msb_FFxDN[45]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n60) );
  DFF_X1 mult_msb_FFxDP_reg_12__1_ ( .D(mult_msb_FFxDN[49]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n43) );
  DFF_X1 mult_msb_FFxDP_reg_13__1_ ( .D(mult_msb_FFxDN[53]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n44) );
  DFF_X1 mult_msb_FFxDP_reg_14__1_ ( .D(mult_msb_FFxDN[57]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n41) );
  DFF_X1 mult_msb_FFxDP_reg_1__2_ ( .D(mult_msb_FFxDN[6]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n88) );
  DFF_X1 mult_msb_FFxDP_reg_2__2_ ( .D(mult_msb_FFxDN[10]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n85) );
  DFF_X1 mult_msb_FFxDP_reg_3__2_ ( .D(mult_msb_FFxDN[14]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n86) );
  DFF_X1 mult_msb_FFxDP_reg_4__2_ ( .D(mult_msb_FFxDN[18]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n71) );
  DFF_X1 mult_msb_FFxDP_reg_6__2_ ( .D(mult_msb_FFxDN[26]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n69) );
  DFF_X1 mult_msb_FFxDP_reg_7__2_ ( .D(mult_msb_FFxDN[30]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n70) );
  DFF_X1 mult_msb_FFxDP_reg_8__2_ ( .D(mult_msb_FFxDN[34]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n53) );
  DFF_X1 mult_msb_FFxDP_reg_9__2_ ( .D(mult_msb_FFxDN[38]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n54) );
  DFF_X1 mult_msb_FFxDP_reg_11__2_ ( .D(mult_msb_FFxDN[46]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n56) );
  DFF_X1 mult_msb_FFxDP_reg_12__2_ ( .D(mult_msb_FFxDN[50]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n39) );
  DFF_X1 mult_msb_FFxDP_reg_13__2_ ( .D(mult_msb_FFxDN[54]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n40) );
  DFF_X1 mult_msb_FFxDP_reg_14__2_ ( .D(mult_msb_FFxDN[58]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n37) );
  DFF_X1 mult_msb_FFxDP_reg_1__0_ ( .D(mult_msb_FFxDN[4]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n96) );
  DFF_X1 mult_msb_FFxDP_reg_2__0_ ( .D(mult_msb_FFxDN[8]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n93) );
  DFF_X1 mult_msb_FFxDP_reg_3__0_ ( .D(mult_msb_FFxDN[12]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n94) );
  DFF_X1 mult_msb_FFxDP_reg_4__0_ ( .D(mult_msb_FFxDN[16]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n79) );
  DFF_X1 mult_msb_FFxDP_reg_6__0_ ( .D(mult_msb_FFxDN[24]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n77) );
  DFF_X1 mult_msb_FFxDP_reg_7__0_ ( .D(mult_msb_FFxDN[28]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n78) );
  DFF_X1 mult_msb_FFxDP_reg_8__0_ ( .D(mult_msb_FFxDN[32]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n61) );
  DFF_X1 mult_msb_FFxDP_reg_9__0_ ( .D(mult_msb_FFxDN[36]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n62) );
  DFF_X1 mult_msb_FFxDP_reg_11__0_ ( .D(mult_msb_FFxDN[44]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n64) );
  DFF_X1 mult_msb_FFxDP_reg_12__0_ ( .D(mult_msb_FFxDN[48]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n47) );
  DFF_X1 mult_msb_FFxDP_reg_13__0_ ( .D(mult_msb_FFxDN[52]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n48) );
  DFF_X1 mult_msb_FFxDP_reg_14__0_ ( .D(mult_msb_FFxDN[56]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n45) );
  DFF_X1 mult_msb_FFxDP_reg_0__3_ ( .D(mult_msb_FFxDN[3]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n83) );
  DFF_X1 mult_msb_FFxDP_reg_5__3_ ( .D(mult_msb_FFxDN[23]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n68) );
  DFF_X1 mult_msb_FFxDP_reg_10__3_ ( .D(mult_msb_FFxDN[43]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n51) );
  DFF_X1 mult_msb_FFxDP_reg_15__3_ ( .D(mult_msb_FFxDN[63]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n34) );
  DFF_X1 mult_msb_FFxDP_reg_0__1_ ( .D(mult_msb_FFxDN[1]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n91) );
  DFF_X1 mult_msb_FFxDP_reg_5__1_ ( .D(mult_msb_FFxDN[21]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n76) );
  DFF_X1 mult_msb_FFxDP_reg_10__1_ ( .D(mult_msb_FFxDN[41]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n59) );
  DFF_X1 mult_msb_FFxDP_reg_15__1_ ( .D(mult_msb_FFxDN[61]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n42) );
  DFF_X1 mult_msb_FFxDP_reg_0__2_ ( .D(mult_msb_FFxDN[2]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n87) );
  DFF_X1 mult_msb_FFxDP_reg_5__2_ ( .D(mult_msb_FFxDN[22]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n72) );
  DFF_X1 mult_msb_FFxDP_reg_10__2_ ( .D(mult_msb_FFxDN[42]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n55) );
  DFF_X1 mult_msb_FFxDP_reg_15__2_ ( .D(mult_msb_FFxDN[62]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n38) );
  DFF_X1 mult_msb_FFxDP_reg_0__0_ ( .D(mult_msb_FFxDN[0]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n95) );
  DFF_X1 mult_msb_FFxDP_reg_5__0_ ( .D(mult_msb_FFxDN[20]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n80) );
  DFF_X1 mult_msb_FFxDP_reg_10__0_ ( .D(mult_msb_FFxDN[40]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n63) );
  DFF_X1 mult_msb_FFxDP_reg_15__0_ ( .D(mult_msb_FFxDN[60]), .CK(ClkxCI), .Q(), 
        .QN(mult_msb_n46) );
  XNOR2_X1 mult_msb_gf4_mul_3_3_U29 ( .A(mult_msb_gf4_mul_3_3_n77), .B(
        mult_msb_gf4_mul_3_3_n76), .ZN(mult_msb_FFxDN[63]) );
  NAND2_X1 mult_msb_gf4_mul_3_3_U28 ( .A1(n119), .A2(Y0_4xDP[15]), .ZN(
        mult_msb_gf4_mul_3_3_n76) );
  XOR2_X1 mult_msb_gf4_mul_3_3_U27 ( .A(mult_msb_gf4_mul_3_3_n75), .B(
        mult_msb_gf4_mul_3_3_n74), .Z(mult_msb_gf4_mul_3_3_n77) );
  XNOR2_X1 mult_msb_gf4_mul_3_3_U26 ( .A(mult_msb_gf4_mul_3_3_n73), .B(
        mult_msb_gf4_mul_3_3_n72), .ZN(mult_msb_FFxDN[62]) );
  NAND2_X1 mult_msb_gf4_mul_3_3_U25 ( .A1(n117), .A2(Y0_4xDP[14]), .ZN(
        mult_msb_gf4_mul_3_3_n72) );
  XOR2_X1 mult_msb_gf4_mul_3_3_U24 ( .A(mult_msb_gf4_mul_3_3_n74), .B(
        mult_msb_gf4_mul_3_3_n71), .Z(mult_msb_gf4_mul_3_3_n73) );
  NOR2_X1 mult_msb_gf4_mul_3_3_U23 ( .A1(mult_msb_gf4_mul_3_3_n70), .A2(
        mult_msb_gf4_mul_3_3_n69), .ZN(mult_msb_gf4_mul_3_3_n74) );
  XNOR2_X1 mult_msb_gf4_mul_3_3_U22 ( .A(n117), .B(n119), .ZN(
        mult_msb_gf4_mul_3_3_n69) );
  XNOR2_X1 mult_msb_gf4_mul_3_3_U21 ( .A(Y0_4xDP[14]), .B(Y0_4xDP[15]), .ZN(
        mult_msb_gf4_mul_3_3_n70) );
  XNOR2_X1 mult_msb_gf4_mul_3_3_U20 ( .A(mult_msb_gf4_mul_3_3_n68), .B(
        mult_msb_gf4_mul_3_3_n67), .ZN(mult_msb_FFxDN[61]) );
  NAND2_X1 mult_msb_gf4_mul_3_3_U19 ( .A1(n115), .A2(Y0_4xDP[13]), .ZN(
        mult_msb_gf4_mul_3_3_n67) );
  XOR2_X1 mult_msb_gf4_mul_3_3_U18 ( .A(mult_msb_gf4_mul_3_3_n75), .B(
        mult_msb_gf4_mul_3_3_n66), .Z(mult_msb_gf4_mul_3_3_n68) );
  XNOR2_X1 mult_msb_gf4_mul_3_3_U17 ( .A(mult_msb_gf4_mul_3_3_n65), .B(
        mult_msb_gf4_mul_3_3_n64), .ZN(mult_msb_gf4_mul_3_3_n75) );
  NAND2_X1 mult_msb_gf4_mul_3_3_U16 ( .A1(mult_msb_gf4_mul_3_3_n63), .A2(
        mult_msb_gf4_mul_3_3_n62), .ZN(mult_msb_gf4_mul_3_3_n64) );
  XNOR2_X1 mult_msb_gf4_mul_3_3_U15 ( .A(mult_msb_gf4_mul_3_3_n61), .B(
        mult_msb_gf4_mul_3_3_n60), .ZN(mult_msb_gf4_mul_3_3_n62) );
  XNOR2_X1 mult_msb_gf4_mul_3_3_U14 ( .A(mult_msb_gf4_mul_3_3_n59), .B(
        mult_msb_gf4_mul_3_3_n58), .ZN(mult_msb_gf4_mul_3_3_n63) );
  XNOR2_X1 mult_msb_gf4_mul_3_3_U13 ( .A(mult_msb_gf4_mul_3_3_n57), .B(
        mult_msb_gf4_mul_3_3_n56), .ZN(mult_msb_FFxDN[60]) );
  NAND2_X1 mult_msb_gf4_mul_3_3_U12 ( .A1(n113), .A2(Y0_4xDP[12]), .ZN(
        mult_msb_gf4_mul_3_3_n56) );
  XOR2_X1 mult_msb_gf4_mul_3_3_U11 ( .A(mult_msb_gf4_mul_3_3_n66), .B(
        mult_msb_gf4_mul_3_3_n71), .Z(mult_msb_gf4_mul_3_3_n57) );
  XNOR2_X1 mult_msb_gf4_mul_3_3_U10 ( .A(mult_msb_gf4_mul_3_3_n55), .B(
        mult_msb_gf4_mul_3_3_n65), .ZN(mult_msb_gf4_mul_3_3_n71) );
  NOR2_X1 mult_msb_gf4_mul_3_3_U9 ( .A1(mult_msb_gf4_mul_3_3_n61), .A2(
        mult_msb_gf4_mul_3_3_n59), .ZN(mult_msb_gf4_mul_3_3_n65) );
  XNOR2_X1 mult_msb_gf4_mul_3_3_U8 ( .A(n113), .B(n117), .ZN(
        mult_msb_gf4_mul_3_3_n59) );
  XNOR2_X1 mult_msb_gf4_mul_3_3_U7 ( .A(Y0_4xDP[12]), .B(Y0_4xDP[14]), .ZN(
        mult_msb_gf4_mul_3_3_n61) );
  NAND2_X1 mult_msb_gf4_mul_3_3_U6 ( .A1(mult_msb_gf4_mul_3_3_n58), .A2(
        mult_msb_gf4_mul_3_3_n60), .ZN(mult_msb_gf4_mul_3_3_n55) );
  XOR2_X1 mult_msb_gf4_mul_3_3_U5 ( .A(Y0_4xDP[13]), .B(Y0_4xDP[15]), .Z(
        mult_msb_gf4_mul_3_3_n60) );
  XOR2_X1 mult_msb_gf4_mul_3_3_U4 ( .A(n115), .B(n119), .Z(
        mult_msb_gf4_mul_3_3_n58) );
  NOR2_X1 mult_msb_gf4_mul_3_3_U3 ( .A1(mult_msb_gf4_mul_3_3_n54), .A2(
        mult_msb_gf4_mul_3_3_n53), .ZN(mult_msb_gf4_mul_3_3_n66) );
  XNOR2_X1 mult_msb_gf4_mul_3_3_U2 ( .A(n113), .B(n115), .ZN(
        mult_msb_gf4_mul_3_3_n53) );
  XNOR2_X1 mult_msb_gf4_mul_3_3_U1 ( .A(Y0_4xDP[12]), .B(Y0_4xDP[13]), .ZN(
        mult_msb_gf4_mul_3_3_n54) );
  XNOR2_X1 mult_msb_gf4_mul_3_2_U29 ( .A(mult_msb_gf4_mul_3_2_n77), .B(
        mult_msb_gf4_mul_3_2_n76), .ZN(mult_msb_Xi_mul_Yj_14__3_) );
  NAND2_X1 mult_msb_gf4_mul_3_2_U28 ( .A1(n119), .A2(Y0_4xDP[11]), .ZN(
        mult_msb_gf4_mul_3_2_n76) );
  XOR2_X1 mult_msb_gf4_mul_3_2_U27 ( .A(mult_msb_gf4_mul_3_2_n75), .B(
        mult_msb_gf4_mul_3_2_n74), .Z(mult_msb_gf4_mul_3_2_n77) );
  XNOR2_X1 mult_msb_gf4_mul_3_2_U26 ( .A(mult_msb_gf4_mul_3_2_n73), .B(
        mult_msb_gf4_mul_3_2_n72), .ZN(mult_msb_Xi_mul_Yj_14__2_) );
  NAND2_X1 mult_msb_gf4_mul_3_2_U25 ( .A1(n117), .A2(Y0_4xDP[10]), .ZN(
        mult_msb_gf4_mul_3_2_n72) );
  XOR2_X1 mult_msb_gf4_mul_3_2_U24 ( .A(mult_msb_gf4_mul_3_2_n74), .B(
        mult_msb_gf4_mul_3_2_n71), .Z(mult_msb_gf4_mul_3_2_n73) );
  NOR2_X1 mult_msb_gf4_mul_3_2_U23 ( .A1(mult_msb_gf4_mul_3_2_n70), .A2(
        mult_msb_gf4_mul_3_2_n69), .ZN(mult_msb_gf4_mul_3_2_n74) );
  XNOR2_X1 mult_msb_gf4_mul_3_2_U22 ( .A(n117), .B(n119), .ZN(
        mult_msb_gf4_mul_3_2_n69) );
  XNOR2_X1 mult_msb_gf4_mul_3_2_U21 ( .A(Y0_4xDP[10]), .B(Y0_4xDP[11]), .ZN(
        mult_msb_gf4_mul_3_2_n70) );
  XNOR2_X1 mult_msb_gf4_mul_3_2_U20 ( .A(mult_msb_gf4_mul_3_2_n68), .B(
        mult_msb_gf4_mul_3_2_n67), .ZN(mult_msb_Xi_mul_Yj_14__1_) );
  NAND2_X1 mult_msb_gf4_mul_3_2_U19 ( .A1(n115), .A2(Y0_4xDP[9]), .ZN(
        mult_msb_gf4_mul_3_2_n67) );
  XOR2_X1 mult_msb_gf4_mul_3_2_U18 ( .A(mult_msb_gf4_mul_3_2_n75), .B(
        mult_msb_gf4_mul_3_2_n66), .Z(mult_msb_gf4_mul_3_2_n68) );
  XNOR2_X1 mult_msb_gf4_mul_3_2_U17 ( .A(mult_msb_gf4_mul_3_2_n65), .B(
        mult_msb_gf4_mul_3_2_n64), .ZN(mult_msb_gf4_mul_3_2_n75) );
  NAND2_X1 mult_msb_gf4_mul_3_2_U16 ( .A1(mult_msb_gf4_mul_3_2_n63), .A2(
        mult_msb_gf4_mul_3_2_n62), .ZN(mult_msb_gf4_mul_3_2_n64) );
  XNOR2_X1 mult_msb_gf4_mul_3_2_U15 ( .A(mult_msb_gf4_mul_3_2_n61), .B(
        mult_msb_gf4_mul_3_2_n60), .ZN(mult_msb_gf4_mul_3_2_n62) );
  XNOR2_X1 mult_msb_gf4_mul_3_2_U14 ( .A(mult_msb_gf4_mul_3_2_n59), .B(
        mult_msb_gf4_mul_3_2_n58), .ZN(mult_msb_gf4_mul_3_2_n63) );
  XNOR2_X1 mult_msb_gf4_mul_3_2_U13 ( .A(mult_msb_gf4_mul_3_2_n57), .B(
        mult_msb_gf4_mul_3_2_n56), .ZN(mult_msb_Xi_mul_Yj_14__0_) );
  NAND2_X1 mult_msb_gf4_mul_3_2_U12 ( .A1(n113), .A2(Y0_4xDP[8]), .ZN(
        mult_msb_gf4_mul_3_2_n56) );
  XOR2_X1 mult_msb_gf4_mul_3_2_U11 ( .A(mult_msb_gf4_mul_3_2_n66), .B(
        mult_msb_gf4_mul_3_2_n71), .Z(mult_msb_gf4_mul_3_2_n57) );
  XNOR2_X1 mult_msb_gf4_mul_3_2_U10 ( .A(mult_msb_gf4_mul_3_2_n55), .B(
        mult_msb_gf4_mul_3_2_n65), .ZN(mult_msb_gf4_mul_3_2_n71) );
  NOR2_X1 mult_msb_gf4_mul_3_2_U9 ( .A1(mult_msb_gf4_mul_3_2_n61), .A2(
        mult_msb_gf4_mul_3_2_n59), .ZN(mult_msb_gf4_mul_3_2_n65) );
  XNOR2_X1 mult_msb_gf4_mul_3_2_U8 ( .A(n113), .B(n117), .ZN(
        mult_msb_gf4_mul_3_2_n59) );
  XNOR2_X1 mult_msb_gf4_mul_3_2_U7 ( .A(Y0_4xDP[8]), .B(Y0_4xDP[10]), .ZN(
        mult_msb_gf4_mul_3_2_n61) );
  NAND2_X1 mult_msb_gf4_mul_3_2_U6 ( .A1(mult_msb_gf4_mul_3_2_n58), .A2(
        mult_msb_gf4_mul_3_2_n60), .ZN(mult_msb_gf4_mul_3_2_n55) );
  XOR2_X1 mult_msb_gf4_mul_3_2_U5 ( .A(Y0_4xDP[9]), .B(Y0_4xDP[11]), .Z(
        mult_msb_gf4_mul_3_2_n60) );
  XOR2_X1 mult_msb_gf4_mul_3_2_U4 ( .A(n115), .B(n119), .Z(
        mult_msb_gf4_mul_3_2_n58) );
  NOR2_X1 mult_msb_gf4_mul_3_2_U3 ( .A1(mult_msb_gf4_mul_3_2_n54), .A2(
        mult_msb_gf4_mul_3_2_n53), .ZN(mult_msb_gf4_mul_3_2_n66) );
  XNOR2_X1 mult_msb_gf4_mul_3_2_U2 ( .A(n113), .B(n115), .ZN(
        mult_msb_gf4_mul_3_2_n53) );
  XNOR2_X1 mult_msb_gf4_mul_3_2_U1 ( .A(Y0_4xDP[8]), .B(Y0_4xDP[9]), .ZN(
        mult_msb_gf4_mul_3_2_n54) );
  XNOR2_X1 mult_msb_gf4_mul_3_1_U29 ( .A(mult_msb_gf4_mul_3_1_n77), .B(
        mult_msb_gf4_mul_3_1_n76), .ZN(mult_msb_Xi_mul_Yj_13__3_) );
  NAND2_X1 mult_msb_gf4_mul_3_1_U28 ( .A1(n119), .A2(Y0_4xDP[7]), .ZN(
        mult_msb_gf4_mul_3_1_n76) );
  XOR2_X1 mult_msb_gf4_mul_3_1_U27 ( .A(mult_msb_gf4_mul_3_1_n75), .B(
        mult_msb_gf4_mul_3_1_n74), .Z(mult_msb_gf4_mul_3_1_n77) );
  XNOR2_X1 mult_msb_gf4_mul_3_1_U26 ( .A(mult_msb_gf4_mul_3_1_n73), .B(
        mult_msb_gf4_mul_3_1_n72), .ZN(mult_msb_Xi_mul_Yj_13__2_) );
  NAND2_X1 mult_msb_gf4_mul_3_1_U25 ( .A1(n117), .A2(Y0_4xDP[6]), .ZN(
        mult_msb_gf4_mul_3_1_n72) );
  XOR2_X1 mult_msb_gf4_mul_3_1_U24 ( .A(mult_msb_gf4_mul_3_1_n74), .B(
        mult_msb_gf4_mul_3_1_n71), .Z(mult_msb_gf4_mul_3_1_n73) );
  NOR2_X1 mult_msb_gf4_mul_3_1_U23 ( .A1(mult_msb_gf4_mul_3_1_n70), .A2(
        mult_msb_gf4_mul_3_1_n69), .ZN(mult_msb_gf4_mul_3_1_n74) );
  XNOR2_X1 mult_msb_gf4_mul_3_1_U22 ( .A(n117), .B(n119), .ZN(
        mult_msb_gf4_mul_3_1_n69) );
  XNOR2_X1 mult_msb_gf4_mul_3_1_U21 ( .A(Y0_4xDP[6]), .B(Y0_4xDP[7]), .ZN(
        mult_msb_gf4_mul_3_1_n70) );
  XNOR2_X1 mult_msb_gf4_mul_3_1_U20 ( .A(mult_msb_gf4_mul_3_1_n68), .B(
        mult_msb_gf4_mul_3_1_n67), .ZN(mult_msb_Xi_mul_Yj_13__1_) );
  NAND2_X1 mult_msb_gf4_mul_3_1_U19 ( .A1(n115), .A2(Y0_4xDP[5]), .ZN(
        mult_msb_gf4_mul_3_1_n67) );
  XOR2_X1 mult_msb_gf4_mul_3_1_U18 ( .A(mult_msb_gf4_mul_3_1_n75), .B(
        mult_msb_gf4_mul_3_1_n66), .Z(mult_msb_gf4_mul_3_1_n68) );
  XNOR2_X1 mult_msb_gf4_mul_3_1_U17 ( .A(mult_msb_gf4_mul_3_1_n65), .B(
        mult_msb_gf4_mul_3_1_n64), .ZN(mult_msb_gf4_mul_3_1_n75) );
  NAND2_X1 mult_msb_gf4_mul_3_1_U16 ( .A1(mult_msb_gf4_mul_3_1_n63), .A2(
        mult_msb_gf4_mul_3_1_n62), .ZN(mult_msb_gf4_mul_3_1_n64) );
  XNOR2_X1 mult_msb_gf4_mul_3_1_U15 ( .A(mult_msb_gf4_mul_3_1_n61), .B(
        mult_msb_gf4_mul_3_1_n60), .ZN(mult_msb_gf4_mul_3_1_n62) );
  XNOR2_X1 mult_msb_gf4_mul_3_1_U14 ( .A(mult_msb_gf4_mul_3_1_n59), .B(
        mult_msb_gf4_mul_3_1_n58), .ZN(mult_msb_gf4_mul_3_1_n63) );
  XNOR2_X1 mult_msb_gf4_mul_3_1_U13 ( .A(mult_msb_gf4_mul_3_1_n57), .B(
        mult_msb_gf4_mul_3_1_n56), .ZN(mult_msb_Xi_mul_Yj_13__0_) );
  NAND2_X1 mult_msb_gf4_mul_3_1_U12 ( .A1(n113), .A2(Y0_4xDP[4]), .ZN(
        mult_msb_gf4_mul_3_1_n56) );
  XOR2_X1 mult_msb_gf4_mul_3_1_U11 ( .A(mult_msb_gf4_mul_3_1_n66), .B(
        mult_msb_gf4_mul_3_1_n71), .Z(mult_msb_gf4_mul_3_1_n57) );
  XNOR2_X1 mult_msb_gf4_mul_3_1_U10 ( .A(mult_msb_gf4_mul_3_1_n55), .B(
        mult_msb_gf4_mul_3_1_n65), .ZN(mult_msb_gf4_mul_3_1_n71) );
  NOR2_X1 mult_msb_gf4_mul_3_1_U9 ( .A1(mult_msb_gf4_mul_3_1_n61), .A2(
        mult_msb_gf4_mul_3_1_n59), .ZN(mult_msb_gf4_mul_3_1_n65) );
  XNOR2_X1 mult_msb_gf4_mul_3_1_U8 ( .A(n113), .B(n117), .ZN(
        mult_msb_gf4_mul_3_1_n59) );
  XNOR2_X1 mult_msb_gf4_mul_3_1_U7 ( .A(Y0_4xDP[4]), .B(Y0_4xDP[6]), .ZN(
        mult_msb_gf4_mul_3_1_n61) );
  NAND2_X1 mult_msb_gf4_mul_3_1_U6 ( .A1(mult_msb_gf4_mul_3_1_n58), .A2(
        mult_msb_gf4_mul_3_1_n60), .ZN(mult_msb_gf4_mul_3_1_n55) );
  XOR2_X1 mult_msb_gf4_mul_3_1_U5 ( .A(Y0_4xDP[5]), .B(Y0_4xDP[7]), .Z(
        mult_msb_gf4_mul_3_1_n60) );
  XOR2_X1 mult_msb_gf4_mul_3_1_U4 ( .A(n115), .B(n119), .Z(
        mult_msb_gf4_mul_3_1_n58) );
  NOR2_X1 mult_msb_gf4_mul_3_1_U3 ( .A1(mult_msb_gf4_mul_3_1_n54), .A2(
        mult_msb_gf4_mul_3_1_n53), .ZN(mult_msb_gf4_mul_3_1_n66) );
  XNOR2_X1 mult_msb_gf4_mul_3_1_U2 ( .A(n113), .B(n115), .ZN(
        mult_msb_gf4_mul_3_1_n53) );
  XNOR2_X1 mult_msb_gf4_mul_3_1_U1 ( .A(Y0_4xDP[4]), .B(Y0_4xDP[5]), .ZN(
        mult_msb_gf4_mul_3_1_n54) );
  XNOR2_X1 mult_msb_gf4_mul_3_0_U29 ( .A(mult_msb_gf4_mul_3_0_n77), .B(
        mult_msb_gf4_mul_3_0_n76), .ZN(mult_msb_Xi_mul_Yj_12__3_) );
  NAND2_X1 mult_msb_gf4_mul_3_0_U28 ( .A1(n119), .A2(Y0_4xDP[3]), .ZN(
        mult_msb_gf4_mul_3_0_n76) );
  XOR2_X1 mult_msb_gf4_mul_3_0_U27 ( .A(mult_msb_gf4_mul_3_0_n75), .B(
        mult_msb_gf4_mul_3_0_n74), .Z(mult_msb_gf4_mul_3_0_n77) );
  XNOR2_X1 mult_msb_gf4_mul_3_0_U26 ( .A(mult_msb_gf4_mul_3_0_n73), .B(
        mult_msb_gf4_mul_3_0_n72), .ZN(mult_msb_Xi_mul_Yj_12__2_) );
  NAND2_X1 mult_msb_gf4_mul_3_0_U25 ( .A1(n117), .A2(Y0_4xDP[2]), .ZN(
        mult_msb_gf4_mul_3_0_n72) );
  XOR2_X1 mult_msb_gf4_mul_3_0_U24 ( .A(mult_msb_gf4_mul_3_0_n74), .B(
        mult_msb_gf4_mul_3_0_n71), .Z(mult_msb_gf4_mul_3_0_n73) );
  NOR2_X1 mult_msb_gf4_mul_3_0_U23 ( .A1(mult_msb_gf4_mul_3_0_n70), .A2(
        mult_msb_gf4_mul_3_0_n69), .ZN(mult_msb_gf4_mul_3_0_n74) );
  XNOR2_X1 mult_msb_gf4_mul_3_0_U22 ( .A(n117), .B(n119), .ZN(
        mult_msb_gf4_mul_3_0_n69) );
  XNOR2_X1 mult_msb_gf4_mul_3_0_U21 ( .A(Y0_4xDP[2]), .B(Y0_4xDP[3]), .ZN(
        mult_msb_gf4_mul_3_0_n70) );
  XNOR2_X1 mult_msb_gf4_mul_3_0_U20 ( .A(mult_msb_gf4_mul_3_0_n68), .B(
        mult_msb_gf4_mul_3_0_n67), .ZN(mult_msb_Xi_mul_Yj_12__1_) );
  NAND2_X1 mult_msb_gf4_mul_3_0_U19 ( .A1(n115), .A2(Y0_4xDP[1]), .ZN(
        mult_msb_gf4_mul_3_0_n67) );
  XOR2_X1 mult_msb_gf4_mul_3_0_U18 ( .A(mult_msb_gf4_mul_3_0_n75), .B(
        mult_msb_gf4_mul_3_0_n66), .Z(mult_msb_gf4_mul_3_0_n68) );
  XNOR2_X1 mult_msb_gf4_mul_3_0_U17 ( .A(mult_msb_gf4_mul_3_0_n65), .B(
        mult_msb_gf4_mul_3_0_n64), .ZN(mult_msb_gf4_mul_3_0_n75) );
  NAND2_X1 mult_msb_gf4_mul_3_0_U16 ( .A1(mult_msb_gf4_mul_3_0_n63), .A2(
        mult_msb_gf4_mul_3_0_n62), .ZN(mult_msb_gf4_mul_3_0_n64) );
  XNOR2_X1 mult_msb_gf4_mul_3_0_U15 ( .A(mult_msb_gf4_mul_3_0_n61), .B(
        mult_msb_gf4_mul_3_0_n60), .ZN(mult_msb_gf4_mul_3_0_n62) );
  XNOR2_X1 mult_msb_gf4_mul_3_0_U14 ( .A(mult_msb_gf4_mul_3_0_n59), .B(
        mult_msb_gf4_mul_3_0_n58), .ZN(mult_msb_gf4_mul_3_0_n63) );
  XNOR2_X1 mult_msb_gf4_mul_3_0_U13 ( .A(mult_msb_gf4_mul_3_0_n57), .B(
        mult_msb_gf4_mul_3_0_n56), .ZN(mult_msb_Xi_mul_Yj_12__0_) );
  NAND2_X1 mult_msb_gf4_mul_3_0_U12 ( .A1(n113), .A2(Y0_4xDP[0]), .ZN(
        mult_msb_gf4_mul_3_0_n56) );
  XOR2_X1 mult_msb_gf4_mul_3_0_U11 ( .A(mult_msb_gf4_mul_3_0_n66), .B(
        mult_msb_gf4_mul_3_0_n71), .Z(mult_msb_gf4_mul_3_0_n57) );
  XNOR2_X1 mult_msb_gf4_mul_3_0_U10 ( .A(mult_msb_gf4_mul_3_0_n55), .B(
        mult_msb_gf4_mul_3_0_n65), .ZN(mult_msb_gf4_mul_3_0_n71) );
  NOR2_X1 mult_msb_gf4_mul_3_0_U9 ( .A1(mult_msb_gf4_mul_3_0_n61), .A2(
        mult_msb_gf4_mul_3_0_n59), .ZN(mult_msb_gf4_mul_3_0_n65) );
  XNOR2_X1 mult_msb_gf4_mul_3_0_U8 ( .A(n113), .B(n117), .ZN(
        mult_msb_gf4_mul_3_0_n59) );
  XNOR2_X1 mult_msb_gf4_mul_3_0_U7 ( .A(Y0_4xDP[0]), .B(Y0_4xDP[2]), .ZN(
        mult_msb_gf4_mul_3_0_n61) );
  NAND2_X1 mult_msb_gf4_mul_3_0_U6 ( .A1(mult_msb_gf4_mul_3_0_n58), .A2(
        mult_msb_gf4_mul_3_0_n60), .ZN(mult_msb_gf4_mul_3_0_n55) );
  XOR2_X1 mult_msb_gf4_mul_3_0_U5 ( .A(Y0_4xDP[1]), .B(Y0_4xDP[3]), .Z(
        mult_msb_gf4_mul_3_0_n60) );
  XOR2_X1 mult_msb_gf4_mul_3_0_U4 ( .A(n115), .B(n119), .Z(
        mult_msb_gf4_mul_3_0_n58) );
  NOR2_X1 mult_msb_gf4_mul_3_0_U3 ( .A1(mult_msb_gf4_mul_3_0_n54), .A2(
        mult_msb_gf4_mul_3_0_n53), .ZN(mult_msb_gf4_mul_3_0_n66) );
  XNOR2_X1 mult_msb_gf4_mul_3_0_U2 ( .A(n113), .B(n115), .ZN(
        mult_msb_gf4_mul_3_0_n53) );
  XNOR2_X1 mult_msb_gf4_mul_3_0_U1 ( .A(Y0_4xDP[0]), .B(Y0_4xDP[1]), .ZN(
        mult_msb_gf4_mul_3_0_n54) );
  XNOR2_X1 mult_msb_gf4_mul_2_3_U29 ( .A(mult_msb_gf4_mul_2_3_n77), .B(
        mult_msb_gf4_mul_2_3_n76), .ZN(mult_msb_Xi_mul_Yj_11__3_) );
  NAND2_X1 mult_msb_gf4_mul_2_3_U28 ( .A1(n111), .A2(Y0_4xDP[15]), .ZN(
        mult_msb_gf4_mul_2_3_n76) );
  XOR2_X1 mult_msb_gf4_mul_2_3_U27 ( .A(mult_msb_gf4_mul_2_3_n75), .B(
        mult_msb_gf4_mul_2_3_n74), .Z(mult_msb_gf4_mul_2_3_n77) );
  XNOR2_X1 mult_msb_gf4_mul_2_3_U26 ( .A(mult_msb_gf4_mul_2_3_n73), .B(
        mult_msb_gf4_mul_2_3_n72), .ZN(mult_msb_Xi_mul_Yj_11__2_) );
  NAND2_X1 mult_msb_gf4_mul_2_3_U25 ( .A1(n109), .A2(Y0_4xDP[14]), .ZN(
        mult_msb_gf4_mul_2_3_n72) );
  XOR2_X1 mult_msb_gf4_mul_2_3_U24 ( .A(mult_msb_gf4_mul_2_3_n74), .B(
        mult_msb_gf4_mul_2_3_n71), .Z(mult_msb_gf4_mul_2_3_n73) );
  NOR2_X1 mult_msb_gf4_mul_2_3_U23 ( .A1(mult_msb_gf4_mul_2_3_n70), .A2(
        mult_msb_gf4_mul_2_3_n69), .ZN(mult_msb_gf4_mul_2_3_n74) );
  XNOR2_X1 mult_msb_gf4_mul_2_3_U22 ( .A(n109), .B(n111), .ZN(
        mult_msb_gf4_mul_2_3_n69) );
  XNOR2_X1 mult_msb_gf4_mul_2_3_U21 ( .A(Y0_4xDP[14]), .B(Y0_4xDP[15]), .ZN(
        mult_msb_gf4_mul_2_3_n70) );
  XNOR2_X1 mult_msb_gf4_mul_2_3_U20 ( .A(mult_msb_gf4_mul_2_3_n68), .B(
        mult_msb_gf4_mul_2_3_n67), .ZN(mult_msb_Xi_mul_Yj_11__1_) );
  NAND2_X1 mult_msb_gf4_mul_2_3_U19 ( .A1(n107), .A2(Y0_4xDP[13]), .ZN(
        mult_msb_gf4_mul_2_3_n67) );
  XOR2_X1 mult_msb_gf4_mul_2_3_U18 ( .A(mult_msb_gf4_mul_2_3_n75), .B(
        mult_msb_gf4_mul_2_3_n66), .Z(mult_msb_gf4_mul_2_3_n68) );
  XNOR2_X1 mult_msb_gf4_mul_2_3_U17 ( .A(mult_msb_gf4_mul_2_3_n65), .B(
        mult_msb_gf4_mul_2_3_n64), .ZN(mult_msb_gf4_mul_2_3_n75) );
  NAND2_X1 mult_msb_gf4_mul_2_3_U16 ( .A1(mult_msb_gf4_mul_2_3_n63), .A2(
        mult_msb_gf4_mul_2_3_n62), .ZN(mult_msb_gf4_mul_2_3_n64) );
  XNOR2_X1 mult_msb_gf4_mul_2_3_U15 ( .A(mult_msb_gf4_mul_2_3_n61), .B(
        mult_msb_gf4_mul_2_3_n60), .ZN(mult_msb_gf4_mul_2_3_n62) );
  XNOR2_X1 mult_msb_gf4_mul_2_3_U14 ( .A(mult_msb_gf4_mul_2_3_n59), .B(
        mult_msb_gf4_mul_2_3_n58), .ZN(mult_msb_gf4_mul_2_3_n63) );
  XNOR2_X1 mult_msb_gf4_mul_2_3_U13 ( .A(mult_msb_gf4_mul_2_3_n57), .B(
        mult_msb_gf4_mul_2_3_n56), .ZN(mult_msb_Xi_mul_Yj_11__0_) );
  NAND2_X1 mult_msb_gf4_mul_2_3_U12 ( .A1(n105), .A2(Y0_4xDP[12]), .ZN(
        mult_msb_gf4_mul_2_3_n56) );
  XOR2_X1 mult_msb_gf4_mul_2_3_U11 ( .A(mult_msb_gf4_mul_2_3_n66), .B(
        mult_msb_gf4_mul_2_3_n71), .Z(mult_msb_gf4_mul_2_3_n57) );
  XNOR2_X1 mult_msb_gf4_mul_2_3_U10 ( .A(mult_msb_gf4_mul_2_3_n55), .B(
        mult_msb_gf4_mul_2_3_n65), .ZN(mult_msb_gf4_mul_2_3_n71) );
  NOR2_X1 mult_msb_gf4_mul_2_3_U9 ( .A1(mult_msb_gf4_mul_2_3_n61), .A2(
        mult_msb_gf4_mul_2_3_n59), .ZN(mult_msb_gf4_mul_2_3_n65) );
  XNOR2_X1 mult_msb_gf4_mul_2_3_U8 ( .A(n105), .B(n109), .ZN(
        mult_msb_gf4_mul_2_3_n59) );
  XNOR2_X1 mult_msb_gf4_mul_2_3_U7 ( .A(Y0_4xDP[12]), .B(Y0_4xDP[14]), .ZN(
        mult_msb_gf4_mul_2_3_n61) );
  NAND2_X1 mult_msb_gf4_mul_2_3_U6 ( .A1(mult_msb_gf4_mul_2_3_n58), .A2(
        mult_msb_gf4_mul_2_3_n60), .ZN(mult_msb_gf4_mul_2_3_n55) );
  XOR2_X1 mult_msb_gf4_mul_2_3_U5 ( .A(Y0_4xDP[13]), .B(Y0_4xDP[15]), .Z(
        mult_msb_gf4_mul_2_3_n60) );
  XOR2_X1 mult_msb_gf4_mul_2_3_U4 ( .A(n107), .B(n111), .Z(
        mult_msb_gf4_mul_2_3_n58) );
  NOR2_X1 mult_msb_gf4_mul_2_3_U3 ( .A1(mult_msb_gf4_mul_2_3_n54), .A2(
        mult_msb_gf4_mul_2_3_n53), .ZN(mult_msb_gf4_mul_2_3_n66) );
  XNOR2_X1 mult_msb_gf4_mul_2_3_U2 ( .A(n105), .B(n107), .ZN(
        mult_msb_gf4_mul_2_3_n53) );
  XNOR2_X1 mult_msb_gf4_mul_2_3_U1 ( .A(Y0_4xDP[12]), .B(Y0_4xDP[13]), .ZN(
        mult_msb_gf4_mul_2_3_n54) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U29 ( .A(mult_msb_gf4_mul_2_2_n77), .B(
        mult_msb_gf4_mul_2_2_n76), .ZN(mult_msb_FFxDN[43]) );
  NAND2_X1 mult_msb_gf4_mul_2_2_U28 ( .A1(n111), .A2(Y0_4xDP[11]), .ZN(
        mult_msb_gf4_mul_2_2_n76) );
  XOR2_X1 mult_msb_gf4_mul_2_2_U27 ( .A(mult_msb_gf4_mul_2_2_n75), .B(
        mult_msb_gf4_mul_2_2_n74), .Z(mult_msb_gf4_mul_2_2_n77) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U26 ( .A(mult_msb_gf4_mul_2_2_n73), .B(
        mult_msb_gf4_mul_2_2_n72), .ZN(mult_msb_FFxDN[42]) );
  NAND2_X1 mult_msb_gf4_mul_2_2_U25 ( .A1(n109), .A2(Y0_4xDP[10]), .ZN(
        mult_msb_gf4_mul_2_2_n72) );
  XOR2_X1 mult_msb_gf4_mul_2_2_U24 ( .A(mult_msb_gf4_mul_2_2_n74), .B(
        mult_msb_gf4_mul_2_2_n71), .Z(mult_msb_gf4_mul_2_2_n73) );
  NOR2_X1 mult_msb_gf4_mul_2_2_U23 ( .A1(mult_msb_gf4_mul_2_2_n70), .A2(
        mult_msb_gf4_mul_2_2_n69), .ZN(mult_msb_gf4_mul_2_2_n74) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U22 ( .A(n109), .B(n111), .ZN(
        mult_msb_gf4_mul_2_2_n69) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U21 ( .A(Y0_4xDP[10]), .B(Y0_4xDP[11]), .ZN(
        mult_msb_gf4_mul_2_2_n70) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U20 ( .A(mult_msb_gf4_mul_2_2_n68), .B(
        mult_msb_gf4_mul_2_2_n67), .ZN(mult_msb_FFxDN[41]) );
  NAND2_X1 mult_msb_gf4_mul_2_2_U19 ( .A1(n107), .A2(Y0_4xDP[9]), .ZN(
        mult_msb_gf4_mul_2_2_n67) );
  XOR2_X1 mult_msb_gf4_mul_2_2_U18 ( .A(mult_msb_gf4_mul_2_2_n75), .B(
        mult_msb_gf4_mul_2_2_n66), .Z(mult_msb_gf4_mul_2_2_n68) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U17 ( .A(mult_msb_gf4_mul_2_2_n65), .B(
        mult_msb_gf4_mul_2_2_n64), .ZN(mult_msb_gf4_mul_2_2_n75) );
  NAND2_X1 mult_msb_gf4_mul_2_2_U16 ( .A1(mult_msb_gf4_mul_2_2_n63), .A2(
        mult_msb_gf4_mul_2_2_n62), .ZN(mult_msb_gf4_mul_2_2_n64) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U15 ( .A(mult_msb_gf4_mul_2_2_n61), .B(
        mult_msb_gf4_mul_2_2_n60), .ZN(mult_msb_gf4_mul_2_2_n62) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U14 ( .A(mult_msb_gf4_mul_2_2_n59), .B(
        mult_msb_gf4_mul_2_2_n58), .ZN(mult_msb_gf4_mul_2_2_n63) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U13 ( .A(mult_msb_gf4_mul_2_2_n57), .B(
        mult_msb_gf4_mul_2_2_n56), .ZN(mult_msb_FFxDN[40]) );
  NAND2_X1 mult_msb_gf4_mul_2_2_U12 ( .A1(n105), .A2(Y0_4xDP[8]), .ZN(
        mult_msb_gf4_mul_2_2_n56) );
  XOR2_X1 mult_msb_gf4_mul_2_2_U11 ( .A(mult_msb_gf4_mul_2_2_n66), .B(
        mult_msb_gf4_mul_2_2_n71), .Z(mult_msb_gf4_mul_2_2_n57) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U10 ( .A(mult_msb_gf4_mul_2_2_n55), .B(
        mult_msb_gf4_mul_2_2_n65), .ZN(mult_msb_gf4_mul_2_2_n71) );
  NOR2_X1 mult_msb_gf4_mul_2_2_U9 ( .A1(mult_msb_gf4_mul_2_2_n61), .A2(
        mult_msb_gf4_mul_2_2_n59), .ZN(mult_msb_gf4_mul_2_2_n65) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U8 ( .A(n105), .B(n109), .ZN(
        mult_msb_gf4_mul_2_2_n59) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U7 ( .A(Y0_4xDP[8]), .B(Y0_4xDP[10]), .ZN(
        mult_msb_gf4_mul_2_2_n61) );
  NAND2_X1 mult_msb_gf4_mul_2_2_U6 ( .A1(mult_msb_gf4_mul_2_2_n58), .A2(
        mult_msb_gf4_mul_2_2_n60), .ZN(mult_msb_gf4_mul_2_2_n55) );
  XOR2_X1 mult_msb_gf4_mul_2_2_U5 ( .A(Y0_4xDP[9]), .B(Y0_4xDP[11]), .Z(
        mult_msb_gf4_mul_2_2_n60) );
  XOR2_X1 mult_msb_gf4_mul_2_2_U4 ( .A(n107), .B(n111), .Z(
        mult_msb_gf4_mul_2_2_n58) );
  NOR2_X1 mult_msb_gf4_mul_2_2_U3 ( .A1(mult_msb_gf4_mul_2_2_n54), .A2(
        mult_msb_gf4_mul_2_2_n53), .ZN(mult_msb_gf4_mul_2_2_n66) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U2 ( .A(n105), .B(n107), .ZN(
        mult_msb_gf4_mul_2_2_n53) );
  XNOR2_X1 mult_msb_gf4_mul_2_2_U1 ( .A(Y0_4xDP[8]), .B(Y0_4xDP[9]), .ZN(
        mult_msb_gf4_mul_2_2_n54) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U29 ( .A(mult_msb_gf4_mul_2_1_n77), .B(
        mult_msb_gf4_mul_2_1_n76), .ZN(mult_msb_Xi_mul_Yj_9__3_) );
  NAND2_X1 mult_msb_gf4_mul_2_1_U28 ( .A1(n111), .A2(Y0_4xDP[7]), .ZN(
        mult_msb_gf4_mul_2_1_n76) );
  XOR2_X1 mult_msb_gf4_mul_2_1_U27 ( .A(mult_msb_gf4_mul_2_1_n75), .B(
        mult_msb_gf4_mul_2_1_n74), .Z(mult_msb_gf4_mul_2_1_n77) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U26 ( .A(mult_msb_gf4_mul_2_1_n73), .B(
        mult_msb_gf4_mul_2_1_n72), .ZN(mult_msb_Xi_mul_Yj_9__2_) );
  NAND2_X1 mult_msb_gf4_mul_2_1_U25 ( .A1(n109), .A2(Y0_4xDP[6]), .ZN(
        mult_msb_gf4_mul_2_1_n72) );
  XOR2_X1 mult_msb_gf4_mul_2_1_U24 ( .A(mult_msb_gf4_mul_2_1_n74), .B(
        mult_msb_gf4_mul_2_1_n71), .Z(mult_msb_gf4_mul_2_1_n73) );
  NOR2_X1 mult_msb_gf4_mul_2_1_U23 ( .A1(mult_msb_gf4_mul_2_1_n70), .A2(
        mult_msb_gf4_mul_2_1_n69), .ZN(mult_msb_gf4_mul_2_1_n74) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U22 ( .A(n109), .B(n111), .ZN(
        mult_msb_gf4_mul_2_1_n69) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U21 ( .A(Y0_4xDP[6]), .B(Y0_4xDP[7]), .ZN(
        mult_msb_gf4_mul_2_1_n70) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U20 ( .A(mult_msb_gf4_mul_2_1_n68), .B(
        mult_msb_gf4_mul_2_1_n67), .ZN(mult_msb_Xi_mul_Yj_9__1_) );
  NAND2_X1 mult_msb_gf4_mul_2_1_U19 ( .A1(n107), .A2(Y0_4xDP[5]), .ZN(
        mult_msb_gf4_mul_2_1_n67) );
  XOR2_X1 mult_msb_gf4_mul_2_1_U18 ( .A(mult_msb_gf4_mul_2_1_n75), .B(
        mult_msb_gf4_mul_2_1_n66), .Z(mult_msb_gf4_mul_2_1_n68) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U17 ( .A(mult_msb_gf4_mul_2_1_n65), .B(
        mult_msb_gf4_mul_2_1_n64), .ZN(mult_msb_gf4_mul_2_1_n75) );
  NAND2_X1 mult_msb_gf4_mul_2_1_U16 ( .A1(mult_msb_gf4_mul_2_1_n63), .A2(
        mult_msb_gf4_mul_2_1_n62), .ZN(mult_msb_gf4_mul_2_1_n64) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U15 ( .A(mult_msb_gf4_mul_2_1_n61), .B(
        mult_msb_gf4_mul_2_1_n60), .ZN(mult_msb_gf4_mul_2_1_n62) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U14 ( .A(mult_msb_gf4_mul_2_1_n59), .B(
        mult_msb_gf4_mul_2_1_n58), .ZN(mult_msb_gf4_mul_2_1_n63) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U13 ( .A(mult_msb_gf4_mul_2_1_n57), .B(
        mult_msb_gf4_mul_2_1_n56), .ZN(mult_msb_Xi_mul_Yj_9__0_) );
  NAND2_X1 mult_msb_gf4_mul_2_1_U12 ( .A1(n105), .A2(Y0_4xDP[4]), .ZN(
        mult_msb_gf4_mul_2_1_n56) );
  XOR2_X1 mult_msb_gf4_mul_2_1_U11 ( .A(mult_msb_gf4_mul_2_1_n66), .B(
        mult_msb_gf4_mul_2_1_n71), .Z(mult_msb_gf4_mul_2_1_n57) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U10 ( .A(mult_msb_gf4_mul_2_1_n55), .B(
        mult_msb_gf4_mul_2_1_n65), .ZN(mult_msb_gf4_mul_2_1_n71) );
  NOR2_X1 mult_msb_gf4_mul_2_1_U9 ( .A1(mult_msb_gf4_mul_2_1_n61), .A2(
        mult_msb_gf4_mul_2_1_n59), .ZN(mult_msb_gf4_mul_2_1_n65) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U8 ( .A(n105), .B(n109), .ZN(
        mult_msb_gf4_mul_2_1_n59) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U7 ( .A(Y0_4xDP[4]), .B(Y0_4xDP[6]), .ZN(
        mult_msb_gf4_mul_2_1_n61) );
  NAND2_X1 mult_msb_gf4_mul_2_1_U6 ( .A1(mult_msb_gf4_mul_2_1_n58), .A2(
        mult_msb_gf4_mul_2_1_n60), .ZN(mult_msb_gf4_mul_2_1_n55) );
  XOR2_X1 mult_msb_gf4_mul_2_1_U5 ( .A(Y0_4xDP[5]), .B(Y0_4xDP[7]), .Z(
        mult_msb_gf4_mul_2_1_n60) );
  XOR2_X1 mult_msb_gf4_mul_2_1_U4 ( .A(n107), .B(n111), .Z(
        mult_msb_gf4_mul_2_1_n58) );
  NOR2_X1 mult_msb_gf4_mul_2_1_U3 ( .A1(mult_msb_gf4_mul_2_1_n54), .A2(
        mult_msb_gf4_mul_2_1_n53), .ZN(mult_msb_gf4_mul_2_1_n66) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U2 ( .A(n105), .B(n107), .ZN(
        mult_msb_gf4_mul_2_1_n53) );
  XNOR2_X1 mult_msb_gf4_mul_2_1_U1 ( .A(Y0_4xDP[4]), .B(Y0_4xDP[5]), .ZN(
        mult_msb_gf4_mul_2_1_n54) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U29 ( .A(mult_msb_gf4_mul_2_0_n77), .B(
        mult_msb_gf4_mul_2_0_n76), .ZN(mult_msb_Xi_mul_Yj_8__3_) );
  NAND2_X1 mult_msb_gf4_mul_2_0_U28 ( .A1(n111), .A2(Y0_4xDP[3]), .ZN(
        mult_msb_gf4_mul_2_0_n76) );
  XOR2_X1 mult_msb_gf4_mul_2_0_U27 ( .A(mult_msb_gf4_mul_2_0_n75), .B(
        mult_msb_gf4_mul_2_0_n74), .Z(mult_msb_gf4_mul_2_0_n77) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U26 ( .A(mult_msb_gf4_mul_2_0_n73), .B(
        mult_msb_gf4_mul_2_0_n72), .ZN(mult_msb_Xi_mul_Yj_8__2_) );
  NAND2_X1 mult_msb_gf4_mul_2_0_U25 ( .A1(n109), .A2(Y0_4xDP[2]), .ZN(
        mult_msb_gf4_mul_2_0_n72) );
  XOR2_X1 mult_msb_gf4_mul_2_0_U24 ( .A(mult_msb_gf4_mul_2_0_n74), .B(
        mult_msb_gf4_mul_2_0_n71), .Z(mult_msb_gf4_mul_2_0_n73) );
  NOR2_X1 mult_msb_gf4_mul_2_0_U23 ( .A1(mult_msb_gf4_mul_2_0_n70), .A2(
        mult_msb_gf4_mul_2_0_n69), .ZN(mult_msb_gf4_mul_2_0_n74) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U22 ( .A(n109), .B(n111), .ZN(
        mult_msb_gf4_mul_2_0_n69) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U21 ( .A(Y0_4xDP[2]), .B(Y0_4xDP[3]), .ZN(
        mult_msb_gf4_mul_2_0_n70) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U20 ( .A(mult_msb_gf4_mul_2_0_n68), .B(
        mult_msb_gf4_mul_2_0_n67), .ZN(mult_msb_Xi_mul_Yj_8__1_) );
  NAND2_X1 mult_msb_gf4_mul_2_0_U19 ( .A1(n107), .A2(Y0_4xDP[1]), .ZN(
        mult_msb_gf4_mul_2_0_n67) );
  XOR2_X1 mult_msb_gf4_mul_2_0_U18 ( .A(mult_msb_gf4_mul_2_0_n75), .B(
        mult_msb_gf4_mul_2_0_n66), .Z(mult_msb_gf4_mul_2_0_n68) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U17 ( .A(mult_msb_gf4_mul_2_0_n65), .B(
        mult_msb_gf4_mul_2_0_n64), .ZN(mult_msb_gf4_mul_2_0_n75) );
  NAND2_X1 mult_msb_gf4_mul_2_0_U16 ( .A1(mult_msb_gf4_mul_2_0_n63), .A2(
        mult_msb_gf4_mul_2_0_n62), .ZN(mult_msb_gf4_mul_2_0_n64) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U15 ( .A(mult_msb_gf4_mul_2_0_n61), .B(
        mult_msb_gf4_mul_2_0_n60), .ZN(mult_msb_gf4_mul_2_0_n62) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U14 ( .A(mult_msb_gf4_mul_2_0_n59), .B(
        mult_msb_gf4_mul_2_0_n58), .ZN(mult_msb_gf4_mul_2_0_n63) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U13 ( .A(mult_msb_gf4_mul_2_0_n57), .B(
        mult_msb_gf4_mul_2_0_n56), .ZN(mult_msb_Xi_mul_Yj_8__0_) );
  NAND2_X1 mult_msb_gf4_mul_2_0_U12 ( .A1(n105), .A2(Y0_4xDP[0]), .ZN(
        mult_msb_gf4_mul_2_0_n56) );
  XOR2_X1 mult_msb_gf4_mul_2_0_U11 ( .A(mult_msb_gf4_mul_2_0_n66), .B(
        mult_msb_gf4_mul_2_0_n71), .Z(mult_msb_gf4_mul_2_0_n57) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U10 ( .A(mult_msb_gf4_mul_2_0_n55), .B(
        mult_msb_gf4_mul_2_0_n65), .ZN(mult_msb_gf4_mul_2_0_n71) );
  NOR2_X1 mult_msb_gf4_mul_2_0_U9 ( .A1(mult_msb_gf4_mul_2_0_n61), .A2(
        mult_msb_gf4_mul_2_0_n59), .ZN(mult_msb_gf4_mul_2_0_n65) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U8 ( .A(n105), .B(n109), .ZN(
        mult_msb_gf4_mul_2_0_n59) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U7 ( .A(Y0_4xDP[0]), .B(Y0_4xDP[2]), .ZN(
        mult_msb_gf4_mul_2_0_n61) );
  NAND2_X1 mult_msb_gf4_mul_2_0_U6 ( .A1(mult_msb_gf4_mul_2_0_n58), .A2(
        mult_msb_gf4_mul_2_0_n60), .ZN(mult_msb_gf4_mul_2_0_n55) );
  XOR2_X1 mult_msb_gf4_mul_2_0_U5 ( .A(Y0_4xDP[1]), .B(Y0_4xDP[3]), .Z(
        mult_msb_gf4_mul_2_0_n60) );
  XOR2_X1 mult_msb_gf4_mul_2_0_U4 ( .A(n107), .B(n111), .Z(
        mult_msb_gf4_mul_2_0_n58) );
  NOR2_X1 mult_msb_gf4_mul_2_0_U3 ( .A1(mult_msb_gf4_mul_2_0_n54), .A2(
        mult_msb_gf4_mul_2_0_n53), .ZN(mult_msb_gf4_mul_2_0_n66) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U2 ( .A(n105), .B(n107), .ZN(
        mult_msb_gf4_mul_2_0_n53) );
  XNOR2_X1 mult_msb_gf4_mul_2_0_U1 ( .A(Y0_4xDP[0]), .B(Y0_4xDP[1]), .ZN(
        mult_msb_gf4_mul_2_0_n54) );
  XNOR2_X1 mult_msb_gf4_mul_1_3_U29 ( .A(mult_msb_gf4_mul_1_3_n77), .B(
        mult_msb_gf4_mul_1_3_n76), .ZN(mult_msb_Xi_mul_Yj_7__3_) );
  NAND2_X1 mult_msb_gf4_mul_1_3_U28 ( .A1(n103), .A2(Y0_4xDP[15]), .ZN(
        mult_msb_gf4_mul_1_3_n76) );
  XOR2_X1 mult_msb_gf4_mul_1_3_U27 ( .A(mult_msb_gf4_mul_1_3_n75), .B(
        mult_msb_gf4_mul_1_3_n74), .Z(mult_msb_gf4_mul_1_3_n77) );
  XNOR2_X1 mult_msb_gf4_mul_1_3_U26 ( .A(mult_msb_gf4_mul_1_3_n73), .B(
        mult_msb_gf4_mul_1_3_n72), .ZN(mult_msb_Xi_mul_Yj_7__2_) );
  NAND2_X1 mult_msb_gf4_mul_1_3_U25 ( .A1(n101), .A2(Y0_4xDP[14]), .ZN(
        mult_msb_gf4_mul_1_3_n72) );
  XOR2_X1 mult_msb_gf4_mul_1_3_U24 ( .A(mult_msb_gf4_mul_1_3_n74), .B(
        mult_msb_gf4_mul_1_3_n71), .Z(mult_msb_gf4_mul_1_3_n73) );
  NOR2_X1 mult_msb_gf4_mul_1_3_U23 ( .A1(mult_msb_gf4_mul_1_3_n70), .A2(
        mult_msb_gf4_mul_1_3_n69), .ZN(mult_msb_gf4_mul_1_3_n74) );
  XNOR2_X1 mult_msb_gf4_mul_1_3_U22 ( .A(n101), .B(n103), .ZN(
        mult_msb_gf4_mul_1_3_n69) );
  XNOR2_X1 mult_msb_gf4_mul_1_3_U21 ( .A(Y0_4xDP[14]), .B(Y0_4xDP[15]), .ZN(
        mult_msb_gf4_mul_1_3_n70) );
  XNOR2_X1 mult_msb_gf4_mul_1_3_U20 ( .A(mult_msb_gf4_mul_1_3_n68), .B(
        mult_msb_gf4_mul_1_3_n67), .ZN(mult_msb_Xi_mul_Yj_7__1_) );
  NAND2_X1 mult_msb_gf4_mul_1_3_U19 ( .A1(n99), .A2(Y0_4xDP[13]), .ZN(
        mult_msb_gf4_mul_1_3_n67) );
  XOR2_X1 mult_msb_gf4_mul_1_3_U18 ( .A(mult_msb_gf4_mul_1_3_n75), .B(
        mult_msb_gf4_mul_1_3_n66), .Z(mult_msb_gf4_mul_1_3_n68) );
  XNOR2_X1 mult_msb_gf4_mul_1_3_U17 ( .A(mult_msb_gf4_mul_1_3_n65), .B(
        mult_msb_gf4_mul_1_3_n64), .ZN(mult_msb_gf4_mul_1_3_n75) );
  NAND2_X1 mult_msb_gf4_mul_1_3_U16 ( .A1(mult_msb_gf4_mul_1_3_n63), .A2(
        mult_msb_gf4_mul_1_3_n62), .ZN(mult_msb_gf4_mul_1_3_n64) );
  XNOR2_X1 mult_msb_gf4_mul_1_3_U15 ( .A(mult_msb_gf4_mul_1_3_n61), .B(
        mult_msb_gf4_mul_1_3_n60), .ZN(mult_msb_gf4_mul_1_3_n62) );
  XNOR2_X1 mult_msb_gf4_mul_1_3_U14 ( .A(mult_msb_gf4_mul_1_3_n59), .B(
        mult_msb_gf4_mul_1_3_n58), .ZN(mult_msb_gf4_mul_1_3_n63) );
  XNOR2_X1 mult_msb_gf4_mul_1_3_U13 ( .A(mult_msb_gf4_mul_1_3_n57), .B(
        mult_msb_gf4_mul_1_3_n56), .ZN(mult_msb_Xi_mul_Yj_7__0_) );
  NAND2_X1 mult_msb_gf4_mul_1_3_U12 ( .A1(n97), .A2(Y0_4xDP[12]), .ZN(
        mult_msb_gf4_mul_1_3_n56) );
  XOR2_X1 mult_msb_gf4_mul_1_3_U11 ( .A(mult_msb_gf4_mul_1_3_n66), .B(
        mult_msb_gf4_mul_1_3_n71), .Z(mult_msb_gf4_mul_1_3_n57) );
  XNOR2_X1 mult_msb_gf4_mul_1_3_U10 ( .A(mult_msb_gf4_mul_1_3_n55), .B(
        mult_msb_gf4_mul_1_3_n65), .ZN(mult_msb_gf4_mul_1_3_n71) );
  NOR2_X1 mult_msb_gf4_mul_1_3_U9 ( .A1(mult_msb_gf4_mul_1_3_n61), .A2(
        mult_msb_gf4_mul_1_3_n59), .ZN(mult_msb_gf4_mul_1_3_n65) );
  XNOR2_X1 mult_msb_gf4_mul_1_3_U8 ( .A(n97), .B(n101), .ZN(
        mult_msb_gf4_mul_1_3_n59) );
  XNOR2_X1 mult_msb_gf4_mul_1_3_U7 ( .A(Y0_4xDP[12]), .B(Y0_4xDP[14]), .ZN(
        mult_msb_gf4_mul_1_3_n61) );
  NAND2_X1 mult_msb_gf4_mul_1_3_U6 ( .A1(mult_msb_gf4_mul_1_3_n58), .A2(
        mult_msb_gf4_mul_1_3_n60), .ZN(mult_msb_gf4_mul_1_3_n55) );
  XOR2_X1 mult_msb_gf4_mul_1_3_U5 ( .A(Y0_4xDP[13]), .B(Y0_4xDP[15]), .Z(
        mult_msb_gf4_mul_1_3_n60) );
  XOR2_X1 mult_msb_gf4_mul_1_3_U4 ( .A(n99), .B(n103), .Z(
        mult_msb_gf4_mul_1_3_n58) );
  NOR2_X1 mult_msb_gf4_mul_1_3_U3 ( .A1(mult_msb_gf4_mul_1_3_n54), .A2(
        mult_msb_gf4_mul_1_3_n53), .ZN(mult_msb_gf4_mul_1_3_n66) );
  XNOR2_X1 mult_msb_gf4_mul_1_3_U2 ( .A(n97), .B(n99), .ZN(
        mult_msb_gf4_mul_1_3_n53) );
  XNOR2_X1 mult_msb_gf4_mul_1_3_U1 ( .A(Y0_4xDP[12]), .B(Y0_4xDP[13]), .ZN(
        mult_msb_gf4_mul_1_3_n54) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U29 ( .A(mult_msb_gf4_mul_1_2_n77), .B(
        mult_msb_gf4_mul_1_2_n76), .ZN(mult_msb_Xi_mul_Yj_6__3_) );
  NAND2_X1 mult_msb_gf4_mul_1_2_U28 ( .A1(n103), .A2(Y0_4xDP[11]), .ZN(
        mult_msb_gf4_mul_1_2_n76) );
  XOR2_X1 mult_msb_gf4_mul_1_2_U27 ( .A(mult_msb_gf4_mul_1_2_n75), .B(
        mult_msb_gf4_mul_1_2_n74), .Z(mult_msb_gf4_mul_1_2_n77) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U26 ( .A(mult_msb_gf4_mul_1_2_n73), .B(
        mult_msb_gf4_mul_1_2_n72), .ZN(mult_msb_Xi_mul_Yj_6__2_) );
  NAND2_X1 mult_msb_gf4_mul_1_2_U25 ( .A1(n101), .A2(Y0_4xDP[10]), .ZN(
        mult_msb_gf4_mul_1_2_n72) );
  XOR2_X1 mult_msb_gf4_mul_1_2_U24 ( .A(mult_msb_gf4_mul_1_2_n74), .B(
        mult_msb_gf4_mul_1_2_n71), .Z(mult_msb_gf4_mul_1_2_n73) );
  NOR2_X1 mult_msb_gf4_mul_1_2_U23 ( .A1(mult_msb_gf4_mul_1_2_n70), .A2(
        mult_msb_gf4_mul_1_2_n69), .ZN(mult_msb_gf4_mul_1_2_n74) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U22 ( .A(n101), .B(n103), .ZN(
        mult_msb_gf4_mul_1_2_n69) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U21 ( .A(Y0_4xDP[10]), .B(Y0_4xDP[11]), .ZN(
        mult_msb_gf4_mul_1_2_n70) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U20 ( .A(mult_msb_gf4_mul_1_2_n68), .B(
        mult_msb_gf4_mul_1_2_n67), .ZN(mult_msb_Xi_mul_Yj_6__1_) );
  NAND2_X1 mult_msb_gf4_mul_1_2_U19 ( .A1(n99), .A2(Y0_4xDP[9]), .ZN(
        mult_msb_gf4_mul_1_2_n67) );
  XOR2_X1 mult_msb_gf4_mul_1_2_U18 ( .A(mult_msb_gf4_mul_1_2_n75), .B(
        mult_msb_gf4_mul_1_2_n66), .Z(mult_msb_gf4_mul_1_2_n68) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U17 ( .A(mult_msb_gf4_mul_1_2_n65), .B(
        mult_msb_gf4_mul_1_2_n64), .ZN(mult_msb_gf4_mul_1_2_n75) );
  NAND2_X1 mult_msb_gf4_mul_1_2_U16 ( .A1(mult_msb_gf4_mul_1_2_n63), .A2(
        mult_msb_gf4_mul_1_2_n62), .ZN(mult_msb_gf4_mul_1_2_n64) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U15 ( .A(mult_msb_gf4_mul_1_2_n61), .B(
        mult_msb_gf4_mul_1_2_n60), .ZN(mult_msb_gf4_mul_1_2_n62) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U14 ( .A(mult_msb_gf4_mul_1_2_n59), .B(
        mult_msb_gf4_mul_1_2_n58), .ZN(mult_msb_gf4_mul_1_2_n63) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U13 ( .A(mult_msb_gf4_mul_1_2_n57), .B(
        mult_msb_gf4_mul_1_2_n56), .ZN(mult_msb_Xi_mul_Yj_6__0_) );
  NAND2_X1 mult_msb_gf4_mul_1_2_U12 ( .A1(n97), .A2(Y0_4xDP[8]), .ZN(
        mult_msb_gf4_mul_1_2_n56) );
  XOR2_X1 mult_msb_gf4_mul_1_2_U11 ( .A(mult_msb_gf4_mul_1_2_n66), .B(
        mult_msb_gf4_mul_1_2_n71), .Z(mult_msb_gf4_mul_1_2_n57) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U10 ( .A(mult_msb_gf4_mul_1_2_n55), .B(
        mult_msb_gf4_mul_1_2_n65), .ZN(mult_msb_gf4_mul_1_2_n71) );
  NOR2_X1 mult_msb_gf4_mul_1_2_U9 ( .A1(mult_msb_gf4_mul_1_2_n61), .A2(
        mult_msb_gf4_mul_1_2_n59), .ZN(mult_msb_gf4_mul_1_2_n65) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U8 ( .A(n97), .B(n101), .ZN(
        mult_msb_gf4_mul_1_2_n59) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U7 ( .A(Y0_4xDP[8]), .B(Y0_4xDP[10]), .ZN(
        mult_msb_gf4_mul_1_2_n61) );
  NAND2_X1 mult_msb_gf4_mul_1_2_U6 ( .A1(mult_msb_gf4_mul_1_2_n58), .A2(
        mult_msb_gf4_mul_1_2_n60), .ZN(mult_msb_gf4_mul_1_2_n55) );
  XOR2_X1 mult_msb_gf4_mul_1_2_U5 ( .A(Y0_4xDP[9]), .B(Y0_4xDP[11]), .Z(
        mult_msb_gf4_mul_1_2_n60) );
  XOR2_X1 mult_msb_gf4_mul_1_2_U4 ( .A(n99), .B(n103), .Z(
        mult_msb_gf4_mul_1_2_n58) );
  NOR2_X1 mult_msb_gf4_mul_1_2_U3 ( .A1(mult_msb_gf4_mul_1_2_n54), .A2(
        mult_msb_gf4_mul_1_2_n53), .ZN(mult_msb_gf4_mul_1_2_n66) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U2 ( .A(n97), .B(n99), .ZN(
        mult_msb_gf4_mul_1_2_n53) );
  XNOR2_X1 mult_msb_gf4_mul_1_2_U1 ( .A(Y0_4xDP[8]), .B(Y0_4xDP[9]), .ZN(
        mult_msb_gf4_mul_1_2_n54) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U29 ( .A(mult_msb_gf4_mul_1_1_n77), .B(
        mult_msb_gf4_mul_1_1_n76), .ZN(mult_msb_FFxDN[23]) );
  NAND2_X1 mult_msb_gf4_mul_1_1_U28 ( .A1(n103), .A2(Y0_4xDP[7]), .ZN(
        mult_msb_gf4_mul_1_1_n76) );
  XOR2_X1 mult_msb_gf4_mul_1_1_U27 ( .A(mult_msb_gf4_mul_1_1_n75), .B(
        mult_msb_gf4_mul_1_1_n74), .Z(mult_msb_gf4_mul_1_1_n77) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U26 ( .A(mult_msb_gf4_mul_1_1_n73), .B(
        mult_msb_gf4_mul_1_1_n72), .ZN(mult_msb_FFxDN[22]) );
  NAND2_X1 mult_msb_gf4_mul_1_1_U25 ( .A1(n101), .A2(Y0_4xDP[6]), .ZN(
        mult_msb_gf4_mul_1_1_n72) );
  XOR2_X1 mult_msb_gf4_mul_1_1_U24 ( .A(mult_msb_gf4_mul_1_1_n74), .B(
        mult_msb_gf4_mul_1_1_n71), .Z(mult_msb_gf4_mul_1_1_n73) );
  NOR2_X1 mult_msb_gf4_mul_1_1_U23 ( .A1(mult_msb_gf4_mul_1_1_n70), .A2(
        mult_msb_gf4_mul_1_1_n69), .ZN(mult_msb_gf4_mul_1_1_n74) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U22 ( .A(n101), .B(n103), .ZN(
        mult_msb_gf4_mul_1_1_n69) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U21 ( .A(Y0_4xDP[6]), .B(Y0_4xDP[7]), .ZN(
        mult_msb_gf4_mul_1_1_n70) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U20 ( .A(mult_msb_gf4_mul_1_1_n68), .B(
        mult_msb_gf4_mul_1_1_n67), .ZN(mult_msb_FFxDN[21]) );
  NAND2_X1 mult_msb_gf4_mul_1_1_U19 ( .A1(n99), .A2(Y0_4xDP[5]), .ZN(
        mult_msb_gf4_mul_1_1_n67) );
  XOR2_X1 mult_msb_gf4_mul_1_1_U18 ( .A(mult_msb_gf4_mul_1_1_n75), .B(
        mult_msb_gf4_mul_1_1_n66), .Z(mult_msb_gf4_mul_1_1_n68) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U17 ( .A(mult_msb_gf4_mul_1_1_n65), .B(
        mult_msb_gf4_mul_1_1_n64), .ZN(mult_msb_gf4_mul_1_1_n75) );
  NAND2_X1 mult_msb_gf4_mul_1_1_U16 ( .A1(mult_msb_gf4_mul_1_1_n63), .A2(
        mult_msb_gf4_mul_1_1_n62), .ZN(mult_msb_gf4_mul_1_1_n64) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U15 ( .A(mult_msb_gf4_mul_1_1_n61), .B(
        mult_msb_gf4_mul_1_1_n60), .ZN(mult_msb_gf4_mul_1_1_n62) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U14 ( .A(mult_msb_gf4_mul_1_1_n59), .B(
        mult_msb_gf4_mul_1_1_n58), .ZN(mult_msb_gf4_mul_1_1_n63) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U13 ( .A(mult_msb_gf4_mul_1_1_n57), .B(
        mult_msb_gf4_mul_1_1_n56), .ZN(mult_msb_FFxDN[20]) );
  NAND2_X1 mult_msb_gf4_mul_1_1_U12 ( .A1(n97), .A2(Y0_4xDP[4]), .ZN(
        mult_msb_gf4_mul_1_1_n56) );
  XOR2_X1 mult_msb_gf4_mul_1_1_U11 ( .A(mult_msb_gf4_mul_1_1_n66), .B(
        mult_msb_gf4_mul_1_1_n71), .Z(mult_msb_gf4_mul_1_1_n57) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U10 ( .A(mult_msb_gf4_mul_1_1_n55), .B(
        mult_msb_gf4_mul_1_1_n65), .ZN(mult_msb_gf4_mul_1_1_n71) );
  NOR2_X1 mult_msb_gf4_mul_1_1_U9 ( .A1(mult_msb_gf4_mul_1_1_n61), .A2(
        mult_msb_gf4_mul_1_1_n59), .ZN(mult_msb_gf4_mul_1_1_n65) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U8 ( .A(n97), .B(n101), .ZN(
        mult_msb_gf4_mul_1_1_n59) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U7 ( .A(Y0_4xDP[4]), .B(Y0_4xDP[6]), .ZN(
        mult_msb_gf4_mul_1_1_n61) );
  NAND2_X1 mult_msb_gf4_mul_1_1_U6 ( .A1(mult_msb_gf4_mul_1_1_n58), .A2(
        mult_msb_gf4_mul_1_1_n60), .ZN(mult_msb_gf4_mul_1_1_n55) );
  XOR2_X1 mult_msb_gf4_mul_1_1_U5 ( .A(Y0_4xDP[5]), .B(Y0_4xDP[7]), .Z(
        mult_msb_gf4_mul_1_1_n60) );
  XOR2_X1 mult_msb_gf4_mul_1_1_U4 ( .A(n99), .B(n103), .Z(
        mult_msb_gf4_mul_1_1_n58) );
  NOR2_X1 mult_msb_gf4_mul_1_1_U3 ( .A1(mult_msb_gf4_mul_1_1_n54), .A2(
        mult_msb_gf4_mul_1_1_n53), .ZN(mult_msb_gf4_mul_1_1_n66) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U2 ( .A(n97), .B(n99), .ZN(
        mult_msb_gf4_mul_1_1_n53) );
  XNOR2_X1 mult_msb_gf4_mul_1_1_U1 ( .A(Y0_4xDP[4]), .B(Y0_4xDP[5]), .ZN(
        mult_msb_gf4_mul_1_1_n54) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U29 ( .A(mult_msb_gf4_mul_1_0_n77), .B(
        mult_msb_gf4_mul_1_0_n76), .ZN(mult_msb_Xi_mul_Yj_4__3_) );
  NAND2_X1 mult_msb_gf4_mul_1_0_U28 ( .A1(n103), .A2(Y0_4xDP[3]), .ZN(
        mult_msb_gf4_mul_1_0_n76) );
  XOR2_X1 mult_msb_gf4_mul_1_0_U27 ( .A(mult_msb_gf4_mul_1_0_n75), .B(
        mult_msb_gf4_mul_1_0_n74), .Z(mult_msb_gf4_mul_1_0_n77) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U26 ( .A(mult_msb_gf4_mul_1_0_n73), .B(
        mult_msb_gf4_mul_1_0_n72), .ZN(mult_msb_Xi_mul_Yj_4__2_) );
  NAND2_X1 mult_msb_gf4_mul_1_0_U25 ( .A1(n101), .A2(Y0_4xDP[2]), .ZN(
        mult_msb_gf4_mul_1_0_n72) );
  XOR2_X1 mult_msb_gf4_mul_1_0_U24 ( .A(mult_msb_gf4_mul_1_0_n74), .B(
        mult_msb_gf4_mul_1_0_n71), .Z(mult_msb_gf4_mul_1_0_n73) );
  NOR2_X1 mult_msb_gf4_mul_1_0_U23 ( .A1(mult_msb_gf4_mul_1_0_n70), .A2(
        mult_msb_gf4_mul_1_0_n69), .ZN(mult_msb_gf4_mul_1_0_n74) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U22 ( .A(n101), .B(n103), .ZN(
        mult_msb_gf4_mul_1_0_n69) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U21 ( .A(Y0_4xDP[2]), .B(Y0_4xDP[3]), .ZN(
        mult_msb_gf4_mul_1_0_n70) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U20 ( .A(mult_msb_gf4_mul_1_0_n68), .B(
        mult_msb_gf4_mul_1_0_n67), .ZN(mult_msb_Xi_mul_Yj_4__1_) );
  NAND2_X1 mult_msb_gf4_mul_1_0_U19 ( .A1(n99), .A2(Y0_4xDP[1]), .ZN(
        mult_msb_gf4_mul_1_0_n67) );
  XOR2_X1 mult_msb_gf4_mul_1_0_U18 ( .A(mult_msb_gf4_mul_1_0_n75), .B(
        mult_msb_gf4_mul_1_0_n66), .Z(mult_msb_gf4_mul_1_0_n68) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U17 ( .A(mult_msb_gf4_mul_1_0_n65), .B(
        mult_msb_gf4_mul_1_0_n64), .ZN(mult_msb_gf4_mul_1_0_n75) );
  NAND2_X1 mult_msb_gf4_mul_1_0_U16 ( .A1(mult_msb_gf4_mul_1_0_n63), .A2(
        mult_msb_gf4_mul_1_0_n62), .ZN(mult_msb_gf4_mul_1_0_n64) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U15 ( .A(mult_msb_gf4_mul_1_0_n61), .B(
        mult_msb_gf4_mul_1_0_n60), .ZN(mult_msb_gf4_mul_1_0_n62) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U14 ( .A(mult_msb_gf4_mul_1_0_n59), .B(
        mult_msb_gf4_mul_1_0_n58), .ZN(mult_msb_gf4_mul_1_0_n63) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U13 ( .A(mult_msb_gf4_mul_1_0_n57), .B(
        mult_msb_gf4_mul_1_0_n56), .ZN(mult_msb_Xi_mul_Yj_4__0_) );
  NAND2_X1 mult_msb_gf4_mul_1_0_U12 ( .A1(n97), .A2(Y0_4xDP[0]), .ZN(
        mult_msb_gf4_mul_1_0_n56) );
  XOR2_X1 mult_msb_gf4_mul_1_0_U11 ( .A(mult_msb_gf4_mul_1_0_n66), .B(
        mult_msb_gf4_mul_1_0_n71), .Z(mult_msb_gf4_mul_1_0_n57) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U10 ( .A(mult_msb_gf4_mul_1_0_n55), .B(
        mult_msb_gf4_mul_1_0_n65), .ZN(mult_msb_gf4_mul_1_0_n71) );
  NOR2_X1 mult_msb_gf4_mul_1_0_U9 ( .A1(mult_msb_gf4_mul_1_0_n61), .A2(
        mult_msb_gf4_mul_1_0_n59), .ZN(mult_msb_gf4_mul_1_0_n65) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U8 ( .A(n97), .B(n101), .ZN(
        mult_msb_gf4_mul_1_0_n59) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U7 ( .A(Y0_4xDP[0]), .B(Y0_4xDP[2]), .ZN(
        mult_msb_gf4_mul_1_0_n61) );
  NAND2_X1 mult_msb_gf4_mul_1_0_U6 ( .A1(mult_msb_gf4_mul_1_0_n58), .A2(
        mult_msb_gf4_mul_1_0_n60), .ZN(mult_msb_gf4_mul_1_0_n55) );
  XOR2_X1 mult_msb_gf4_mul_1_0_U5 ( .A(Y0_4xDP[1]), .B(Y0_4xDP[3]), .Z(
        mult_msb_gf4_mul_1_0_n60) );
  XOR2_X1 mult_msb_gf4_mul_1_0_U4 ( .A(n99), .B(n103), .Z(
        mult_msb_gf4_mul_1_0_n58) );
  NOR2_X1 mult_msb_gf4_mul_1_0_U3 ( .A1(mult_msb_gf4_mul_1_0_n54), .A2(
        mult_msb_gf4_mul_1_0_n53), .ZN(mult_msb_gf4_mul_1_0_n66) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U2 ( .A(n97), .B(n99), .ZN(
        mult_msb_gf4_mul_1_0_n53) );
  XNOR2_X1 mult_msb_gf4_mul_1_0_U1 ( .A(Y0_4xDP[0]), .B(Y0_4xDP[1]), .ZN(
        mult_msb_gf4_mul_1_0_n54) );
  XNOR2_X1 mult_msb_gf4_mul_0_3_U29 ( .A(mult_msb_gf4_mul_0_3_n77), .B(
        mult_msb_gf4_mul_0_3_n76), .ZN(mult_msb_Xi_mul_Yj_3__3_) );
  NAND2_X1 mult_msb_gf4_mul_0_3_U28 ( .A1(n95), .A2(Y0_4xDP[15]), .ZN(
        mult_msb_gf4_mul_0_3_n76) );
  XOR2_X1 mult_msb_gf4_mul_0_3_U27 ( .A(mult_msb_gf4_mul_0_3_n75), .B(
        mult_msb_gf4_mul_0_3_n74), .Z(mult_msb_gf4_mul_0_3_n77) );
  XNOR2_X1 mult_msb_gf4_mul_0_3_U26 ( .A(mult_msb_gf4_mul_0_3_n73), .B(
        mult_msb_gf4_mul_0_3_n72), .ZN(mult_msb_Xi_mul_Yj_3__2_) );
  NAND2_X1 mult_msb_gf4_mul_0_3_U25 ( .A1(n93), .A2(Y0_4xDP[14]), .ZN(
        mult_msb_gf4_mul_0_3_n72) );
  XOR2_X1 mult_msb_gf4_mul_0_3_U24 ( .A(mult_msb_gf4_mul_0_3_n74), .B(
        mult_msb_gf4_mul_0_3_n71), .Z(mult_msb_gf4_mul_0_3_n73) );
  NOR2_X1 mult_msb_gf4_mul_0_3_U23 ( .A1(mult_msb_gf4_mul_0_3_n70), .A2(
        mult_msb_gf4_mul_0_3_n69), .ZN(mult_msb_gf4_mul_0_3_n74) );
  XNOR2_X1 mult_msb_gf4_mul_0_3_U22 ( .A(n93), .B(n95), .ZN(
        mult_msb_gf4_mul_0_3_n69) );
  XNOR2_X1 mult_msb_gf4_mul_0_3_U21 ( .A(Y0_4xDP[14]), .B(Y0_4xDP[15]), .ZN(
        mult_msb_gf4_mul_0_3_n70) );
  XNOR2_X1 mult_msb_gf4_mul_0_3_U20 ( .A(mult_msb_gf4_mul_0_3_n68), .B(
        mult_msb_gf4_mul_0_3_n67), .ZN(mult_msb_Xi_mul_Yj_3__1_) );
  NAND2_X1 mult_msb_gf4_mul_0_3_U19 ( .A1(n91), .A2(Y0_4xDP[13]), .ZN(
        mult_msb_gf4_mul_0_3_n67) );
  XOR2_X1 mult_msb_gf4_mul_0_3_U18 ( .A(mult_msb_gf4_mul_0_3_n75), .B(
        mult_msb_gf4_mul_0_3_n66), .Z(mult_msb_gf4_mul_0_3_n68) );
  XNOR2_X1 mult_msb_gf4_mul_0_3_U17 ( .A(mult_msb_gf4_mul_0_3_n65), .B(
        mult_msb_gf4_mul_0_3_n64), .ZN(mult_msb_gf4_mul_0_3_n75) );
  NAND2_X1 mult_msb_gf4_mul_0_3_U16 ( .A1(mult_msb_gf4_mul_0_3_n63), .A2(
        mult_msb_gf4_mul_0_3_n62), .ZN(mult_msb_gf4_mul_0_3_n64) );
  XNOR2_X1 mult_msb_gf4_mul_0_3_U15 ( .A(mult_msb_gf4_mul_0_3_n61), .B(
        mult_msb_gf4_mul_0_3_n60), .ZN(mult_msb_gf4_mul_0_3_n62) );
  XNOR2_X1 mult_msb_gf4_mul_0_3_U14 ( .A(mult_msb_gf4_mul_0_3_n59), .B(
        mult_msb_gf4_mul_0_3_n58), .ZN(mult_msb_gf4_mul_0_3_n63) );
  XNOR2_X1 mult_msb_gf4_mul_0_3_U13 ( .A(mult_msb_gf4_mul_0_3_n57), .B(
        mult_msb_gf4_mul_0_3_n56), .ZN(mult_msb_Xi_mul_Yj_3__0_) );
  NAND2_X1 mult_msb_gf4_mul_0_3_U12 ( .A1(n89), .A2(Y0_4xDP[12]), .ZN(
        mult_msb_gf4_mul_0_3_n56) );
  XOR2_X1 mult_msb_gf4_mul_0_3_U11 ( .A(mult_msb_gf4_mul_0_3_n66), .B(
        mult_msb_gf4_mul_0_3_n71), .Z(mult_msb_gf4_mul_0_3_n57) );
  XNOR2_X1 mult_msb_gf4_mul_0_3_U10 ( .A(mult_msb_gf4_mul_0_3_n55), .B(
        mult_msb_gf4_mul_0_3_n65), .ZN(mult_msb_gf4_mul_0_3_n71) );
  NOR2_X1 mult_msb_gf4_mul_0_3_U9 ( .A1(mult_msb_gf4_mul_0_3_n61), .A2(
        mult_msb_gf4_mul_0_3_n59), .ZN(mult_msb_gf4_mul_0_3_n65) );
  XNOR2_X1 mult_msb_gf4_mul_0_3_U8 ( .A(n89), .B(n93), .ZN(
        mult_msb_gf4_mul_0_3_n59) );
  XNOR2_X1 mult_msb_gf4_mul_0_3_U7 ( .A(Y0_4xDP[12]), .B(Y0_4xDP[14]), .ZN(
        mult_msb_gf4_mul_0_3_n61) );
  NAND2_X1 mult_msb_gf4_mul_0_3_U6 ( .A1(mult_msb_gf4_mul_0_3_n58), .A2(
        mult_msb_gf4_mul_0_3_n60), .ZN(mult_msb_gf4_mul_0_3_n55) );
  XOR2_X1 mult_msb_gf4_mul_0_3_U5 ( .A(Y0_4xDP[13]), .B(Y0_4xDP[15]), .Z(
        mult_msb_gf4_mul_0_3_n60) );
  XOR2_X1 mult_msb_gf4_mul_0_3_U4 ( .A(n91), .B(n95), .Z(
        mult_msb_gf4_mul_0_3_n58) );
  NOR2_X1 mult_msb_gf4_mul_0_3_U3 ( .A1(mult_msb_gf4_mul_0_3_n54), .A2(
        mult_msb_gf4_mul_0_3_n53), .ZN(mult_msb_gf4_mul_0_3_n66) );
  XNOR2_X1 mult_msb_gf4_mul_0_3_U2 ( .A(n89), .B(n91), .ZN(
        mult_msb_gf4_mul_0_3_n53) );
  XNOR2_X1 mult_msb_gf4_mul_0_3_U1 ( .A(Y0_4xDP[12]), .B(Y0_4xDP[13]), .ZN(
        mult_msb_gf4_mul_0_3_n54) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U29 ( .A(mult_msb_gf4_mul_0_2_n77), .B(
        mult_msb_gf4_mul_0_2_n76), .ZN(mult_msb_Xi_mul_Yj_2__3_) );
  NAND2_X1 mult_msb_gf4_mul_0_2_U28 ( .A1(n95), .A2(Y0_4xDP[11]), .ZN(
        mult_msb_gf4_mul_0_2_n76) );
  XOR2_X1 mult_msb_gf4_mul_0_2_U27 ( .A(mult_msb_gf4_mul_0_2_n75), .B(
        mult_msb_gf4_mul_0_2_n74), .Z(mult_msb_gf4_mul_0_2_n77) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U26 ( .A(mult_msb_gf4_mul_0_2_n73), .B(
        mult_msb_gf4_mul_0_2_n72), .ZN(mult_msb_Xi_mul_Yj_2__2_) );
  NAND2_X1 mult_msb_gf4_mul_0_2_U25 ( .A1(n93), .A2(Y0_4xDP[10]), .ZN(
        mult_msb_gf4_mul_0_2_n72) );
  XOR2_X1 mult_msb_gf4_mul_0_2_U24 ( .A(mult_msb_gf4_mul_0_2_n74), .B(
        mult_msb_gf4_mul_0_2_n71), .Z(mult_msb_gf4_mul_0_2_n73) );
  NOR2_X1 mult_msb_gf4_mul_0_2_U23 ( .A1(mult_msb_gf4_mul_0_2_n70), .A2(
        mult_msb_gf4_mul_0_2_n69), .ZN(mult_msb_gf4_mul_0_2_n74) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U22 ( .A(n93), .B(n95), .ZN(
        mult_msb_gf4_mul_0_2_n69) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U21 ( .A(Y0_4xDP[10]), .B(Y0_4xDP[11]), .ZN(
        mult_msb_gf4_mul_0_2_n70) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U20 ( .A(mult_msb_gf4_mul_0_2_n68), .B(
        mult_msb_gf4_mul_0_2_n67), .ZN(mult_msb_Xi_mul_Yj_2__1_) );
  NAND2_X1 mult_msb_gf4_mul_0_2_U19 ( .A1(n91), .A2(Y0_4xDP[9]), .ZN(
        mult_msb_gf4_mul_0_2_n67) );
  XOR2_X1 mult_msb_gf4_mul_0_2_U18 ( .A(mult_msb_gf4_mul_0_2_n75), .B(
        mult_msb_gf4_mul_0_2_n66), .Z(mult_msb_gf4_mul_0_2_n68) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U17 ( .A(mult_msb_gf4_mul_0_2_n65), .B(
        mult_msb_gf4_mul_0_2_n64), .ZN(mult_msb_gf4_mul_0_2_n75) );
  NAND2_X1 mult_msb_gf4_mul_0_2_U16 ( .A1(mult_msb_gf4_mul_0_2_n63), .A2(
        mult_msb_gf4_mul_0_2_n62), .ZN(mult_msb_gf4_mul_0_2_n64) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U15 ( .A(mult_msb_gf4_mul_0_2_n61), .B(
        mult_msb_gf4_mul_0_2_n60), .ZN(mult_msb_gf4_mul_0_2_n62) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U14 ( .A(mult_msb_gf4_mul_0_2_n59), .B(
        mult_msb_gf4_mul_0_2_n58), .ZN(mult_msb_gf4_mul_0_2_n63) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U13 ( .A(mult_msb_gf4_mul_0_2_n57), .B(
        mult_msb_gf4_mul_0_2_n56), .ZN(mult_msb_Xi_mul_Yj_2__0_) );
  NAND2_X1 mult_msb_gf4_mul_0_2_U12 ( .A1(n89), .A2(Y0_4xDP[8]), .ZN(
        mult_msb_gf4_mul_0_2_n56) );
  XOR2_X1 mult_msb_gf4_mul_0_2_U11 ( .A(mult_msb_gf4_mul_0_2_n66), .B(
        mult_msb_gf4_mul_0_2_n71), .Z(mult_msb_gf4_mul_0_2_n57) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U10 ( .A(mult_msb_gf4_mul_0_2_n55), .B(
        mult_msb_gf4_mul_0_2_n65), .ZN(mult_msb_gf4_mul_0_2_n71) );
  NOR2_X1 mult_msb_gf4_mul_0_2_U9 ( .A1(mult_msb_gf4_mul_0_2_n61), .A2(
        mult_msb_gf4_mul_0_2_n59), .ZN(mult_msb_gf4_mul_0_2_n65) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U8 ( .A(n89), .B(n93), .ZN(
        mult_msb_gf4_mul_0_2_n59) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U7 ( .A(Y0_4xDP[8]), .B(Y0_4xDP[10]), .ZN(
        mult_msb_gf4_mul_0_2_n61) );
  NAND2_X1 mult_msb_gf4_mul_0_2_U6 ( .A1(mult_msb_gf4_mul_0_2_n58), .A2(
        mult_msb_gf4_mul_0_2_n60), .ZN(mult_msb_gf4_mul_0_2_n55) );
  XOR2_X1 mult_msb_gf4_mul_0_2_U5 ( .A(Y0_4xDP[9]), .B(Y0_4xDP[11]), .Z(
        mult_msb_gf4_mul_0_2_n60) );
  XOR2_X1 mult_msb_gf4_mul_0_2_U4 ( .A(n91), .B(n95), .Z(
        mult_msb_gf4_mul_0_2_n58) );
  NOR2_X1 mult_msb_gf4_mul_0_2_U3 ( .A1(mult_msb_gf4_mul_0_2_n54), .A2(
        mult_msb_gf4_mul_0_2_n53), .ZN(mult_msb_gf4_mul_0_2_n66) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U2 ( .A(n89), .B(n91), .ZN(
        mult_msb_gf4_mul_0_2_n53) );
  XNOR2_X1 mult_msb_gf4_mul_0_2_U1 ( .A(Y0_4xDP[8]), .B(Y0_4xDP[9]), .ZN(
        mult_msb_gf4_mul_0_2_n54) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U29 ( .A(mult_msb_gf4_mul_0_1_n77), .B(
        mult_msb_gf4_mul_0_1_n76), .ZN(mult_msb_Xi_mul_Yj_1__3_) );
  NAND2_X1 mult_msb_gf4_mul_0_1_U28 ( .A1(n95), .A2(Y0_4xDP[7]), .ZN(
        mult_msb_gf4_mul_0_1_n76) );
  XOR2_X1 mult_msb_gf4_mul_0_1_U27 ( .A(mult_msb_gf4_mul_0_1_n75), .B(
        mult_msb_gf4_mul_0_1_n74), .Z(mult_msb_gf4_mul_0_1_n77) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U26 ( .A(mult_msb_gf4_mul_0_1_n73), .B(
        mult_msb_gf4_mul_0_1_n72), .ZN(mult_msb_Xi_mul_Yj_1__2_) );
  NAND2_X1 mult_msb_gf4_mul_0_1_U25 ( .A1(n93), .A2(Y0_4xDP[6]), .ZN(
        mult_msb_gf4_mul_0_1_n72) );
  XOR2_X1 mult_msb_gf4_mul_0_1_U24 ( .A(mult_msb_gf4_mul_0_1_n74), .B(
        mult_msb_gf4_mul_0_1_n71), .Z(mult_msb_gf4_mul_0_1_n73) );
  NOR2_X1 mult_msb_gf4_mul_0_1_U23 ( .A1(mult_msb_gf4_mul_0_1_n70), .A2(
        mult_msb_gf4_mul_0_1_n69), .ZN(mult_msb_gf4_mul_0_1_n74) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U22 ( .A(n93), .B(n95), .ZN(
        mult_msb_gf4_mul_0_1_n69) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U21 ( .A(Y0_4xDP[6]), .B(Y0_4xDP[7]), .ZN(
        mult_msb_gf4_mul_0_1_n70) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U20 ( .A(mult_msb_gf4_mul_0_1_n68), .B(
        mult_msb_gf4_mul_0_1_n67), .ZN(mult_msb_Xi_mul_Yj_1__1_) );
  NAND2_X1 mult_msb_gf4_mul_0_1_U19 ( .A1(n91), .A2(Y0_4xDP[5]), .ZN(
        mult_msb_gf4_mul_0_1_n67) );
  XOR2_X1 mult_msb_gf4_mul_0_1_U18 ( .A(mult_msb_gf4_mul_0_1_n75), .B(
        mult_msb_gf4_mul_0_1_n66), .Z(mult_msb_gf4_mul_0_1_n68) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U17 ( .A(mult_msb_gf4_mul_0_1_n65), .B(
        mult_msb_gf4_mul_0_1_n64), .ZN(mult_msb_gf4_mul_0_1_n75) );
  NAND2_X1 mult_msb_gf4_mul_0_1_U16 ( .A1(mult_msb_gf4_mul_0_1_n63), .A2(
        mult_msb_gf4_mul_0_1_n62), .ZN(mult_msb_gf4_mul_0_1_n64) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U15 ( .A(mult_msb_gf4_mul_0_1_n61), .B(
        mult_msb_gf4_mul_0_1_n60), .ZN(mult_msb_gf4_mul_0_1_n62) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U14 ( .A(mult_msb_gf4_mul_0_1_n59), .B(
        mult_msb_gf4_mul_0_1_n58), .ZN(mult_msb_gf4_mul_0_1_n63) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U13 ( .A(mult_msb_gf4_mul_0_1_n57), .B(
        mult_msb_gf4_mul_0_1_n56), .ZN(mult_msb_Xi_mul_Yj_1__0_) );
  NAND2_X1 mult_msb_gf4_mul_0_1_U12 ( .A1(n89), .A2(Y0_4xDP[4]), .ZN(
        mult_msb_gf4_mul_0_1_n56) );
  XOR2_X1 mult_msb_gf4_mul_0_1_U11 ( .A(mult_msb_gf4_mul_0_1_n66), .B(
        mult_msb_gf4_mul_0_1_n71), .Z(mult_msb_gf4_mul_0_1_n57) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U10 ( .A(mult_msb_gf4_mul_0_1_n55), .B(
        mult_msb_gf4_mul_0_1_n65), .ZN(mult_msb_gf4_mul_0_1_n71) );
  NOR2_X1 mult_msb_gf4_mul_0_1_U9 ( .A1(mult_msb_gf4_mul_0_1_n61), .A2(
        mult_msb_gf4_mul_0_1_n59), .ZN(mult_msb_gf4_mul_0_1_n65) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U8 ( .A(n89), .B(n93), .ZN(
        mult_msb_gf4_mul_0_1_n59) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U7 ( .A(Y0_4xDP[4]), .B(Y0_4xDP[6]), .ZN(
        mult_msb_gf4_mul_0_1_n61) );
  NAND2_X1 mult_msb_gf4_mul_0_1_U6 ( .A1(mult_msb_gf4_mul_0_1_n58), .A2(
        mult_msb_gf4_mul_0_1_n60), .ZN(mult_msb_gf4_mul_0_1_n55) );
  XOR2_X1 mult_msb_gf4_mul_0_1_U5 ( .A(Y0_4xDP[5]), .B(Y0_4xDP[7]), .Z(
        mult_msb_gf4_mul_0_1_n60) );
  XOR2_X1 mult_msb_gf4_mul_0_1_U4 ( .A(n91), .B(n95), .Z(
        mult_msb_gf4_mul_0_1_n58) );
  NOR2_X1 mult_msb_gf4_mul_0_1_U3 ( .A1(mult_msb_gf4_mul_0_1_n54), .A2(
        mult_msb_gf4_mul_0_1_n53), .ZN(mult_msb_gf4_mul_0_1_n66) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U2 ( .A(n89), .B(n91), .ZN(
        mult_msb_gf4_mul_0_1_n53) );
  XNOR2_X1 mult_msb_gf4_mul_0_1_U1 ( .A(Y0_4xDP[4]), .B(Y0_4xDP[5]), .ZN(
        mult_msb_gf4_mul_0_1_n54) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U29 ( .A(mult_msb_gf4_mul_0_0_n77), .B(
        mult_msb_gf4_mul_0_0_n76), .ZN(mult_msb_FFxDN[3]) );
  NAND2_X1 mult_msb_gf4_mul_0_0_U28 ( .A1(n95), .A2(Y0_4xDP[3]), .ZN(
        mult_msb_gf4_mul_0_0_n76) );
  XOR2_X1 mult_msb_gf4_mul_0_0_U27 ( .A(mult_msb_gf4_mul_0_0_n75), .B(
        mult_msb_gf4_mul_0_0_n74), .Z(mult_msb_gf4_mul_0_0_n77) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U26 ( .A(mult_msb_gf4_mul_0_0_n73), .B(
        mult_msb_gf4_mul_0_0_n72), .ZN(mult_msb_FFxDN[2]) );
  NAND2_X1 mult_msb_gf4_mul_0_0_U25 ( .A1(n93), .A2(Y0_4xDP[2]), .ZN(
        mult_msb_gf4_mul_0_0_n72) );
  XOR2_X1 mult_msb_gf4_mul_0_0_U24 ( .A(mult_msb_gf4_mul_0_0_n74), .B(
        mult_msb_gf4_mul_0_0_n71), .Z(mult_msb_gf4_mul_0_0_n73) );
  NOR2_X1 mult_msb_gf4_mul_0_0_U23 ( .A1(mult_msb_gf4_mul_0_0_n70), .A2(
        mult_msb_gf4_mul_0_0_n69), .ZN(mult_msb_gf4_mul_0_0_n74) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U22 ( .A(n93), .B(n95), .ZN(
        mult_msb_gf4_mul_0_0_n69) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U21 ( .A(Y0_4xDP[2]), .B(Y0_4xDP[3]), .ZN(
        mult_msb_gf4_mul_0_0_n70) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U20 ( .A(mult_msb_gf4_mul_0_0_n68), .B(
        mult_msb_gf4_mul_0_0_n67), .ZN(mult_msb_FFxDN[1]) );
  NAND2_X1 mult_msb_gf4_mul_0_0_U19 ( .A1(n91), .A2(Y0_4xDP[1]), .ZN(
        mult_msb_gf4_mul_0_0_n67) );
  XOR2_X1 mult_msb_gf4_mul_0_0_U18 ( .A(mult_msb_gf4_mul_0_0_n75), .B(
        mult_msb_gf4_mul_0_0_n66), .Z(mult_msb_gf4_mul_0_0_n68) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U17 ( .A(mult_msb_gf4_mul_0_0_n65), .B(
        mult_msb_gf4_mul_0_0_n64), .ZN(mult_msb_gf4_mul_0_0_n75) );
  NAND2_X1 mult_msb_gf4_mul_0_0_U16 ( .A1(mult_msb_gf4_mul_0_0_n63), .A2(
        mult_msb_gf4_mul_0_0_n62), .ZN(mult_msb_gf4_mul_0_0_n64) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U15 ( .A(mult_msb_gf4_mul_0_0_n61), .B(
        mult_msb_gf4_mul_0_0_n60), .ZN(mult_msb_gf4_mul_0_0_n62) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U14 ( .A(mult_msb_gf4_mul_0_0_n59), .B(
        mult_msb_gf4_mul_0_0_n58), .ZN(mult_msb_gf4_mul_0_0_n63) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U13 ( .A(mult_msb_gf4_mul_0_0_n57), .B(
        mult_msb_gf4_mul_0_0_n56), .ZN(mult_msb_FFxDN[0]) );
  NAND2_X1 mult_msb_gf4_mul_0_0_U12 ( .A1(n89), .A2(Y0_4xDP[0]), .ZN(
        mult_msb_gf4_mul_0_0_n56) );
  XOR2_X1 mult_msb_gf4_mul_0_0_U11 ( .A(mult_msb_gf4_mul_0_0_n66), .B(
        mult_msb_gf4_mul_0_0_n71), .Z(mult_msb_gf4_mul_0_0_n57) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U10 ( .A(mult_msb_gf4_mul_0_0_n55), .B(
        mult_msb_gf4_mul_0_0_n65), .ZN(mult_msb_gf4_mul_0_0_n71) );
  NOR2_X1 mult_msb_gf4_mul_0_0_U9 ( .A1(mult_msb_gf4_mul_0_0_n61), .A2(
        mult_msb_gf4_mul_0_0_n59), .ZN(mult_msb_gf4_mul_0_0_n65) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U8 ( .A(n89), .B(n93), .ZN(
        mult_msb_gf4_mul_0_0_n59) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U7 ( .A(Y0_4xDP[0]), .B(Y0_4xDP[2]), .ZN(
        mult_msb_gf4_mul_0_0_n61) );
  NAND2_X1 mult_msb_gf4_mul_0_0_U6 ( .A1(mult_msb_gf4_mul_0_0_n58), .A2(
        mult_msb_gf4_mul_0_0_n60), .ZN(mult_msb_gf4_mul_0_0_n55) );
  XOR2_X1 mult_msb_gf4_mul_0_0_U5 ( .A(Y0_4xDP[1]), .B(Y0_4xDP[3]), .Z(
        mult_msb_gf4_mul_0_0_n60) );
  XOR2_X1 mult_msb_gf4_mul_0_0_U4 ( .A(n91), .B(n95), .Z(
        mult_msb_gf4_mul_0_0_n58) );
  NOR2_X1 mult_msb_gf4_mul_0_0_U3 ( .A1(mult_msb_gf4_mul_0_0_n54), .A2(
        mult_msb_gf4_mul_0_0_n53), .ZN(mult_msb_gf4_mul_0_0_n66) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U2 ( .A(n89), .B(n91), .ZN(
        mult_msb_gf4_mul_0_0_n53) );
  XNOR2_X1 mult_msb_gf4_mul_0_0_U1 ( .A(Y0_4xDP[0]), .B(Y0_4xDP[1]), .ZN(
        mult_msb_gf4_mul_0_0_n54) );
  XNOR2_X1 mult_lsb_U98 ( .A(mult_lsb_n128), .B(mult_lsb_n127), .ZN(
        InvUnmappedxD[27]) );
  XNOR2_X1 mult_lsb_U97 ( .A(mult_lsb_n34), .B(mult_lsb_n33), .ZN(
        mult_lsb_n127) );
  XOR2_X1 mult_lsb_U96 ( .A(mult_lsb_n36), .B(mult_lsb_n35), .Z(mult_lsb_n128)
         );
  XNOR2_X1 mult_lsb_U95 ( .A(mult_lsb_n126), .B(mult_lsb_n125), .ZN(
        InvUnmappedxD[26]) );
  XNOR2_X1 mult_lsb_U94 ( .A(mult_lsb_n38), .B(mult_lsb_n37), .ZN(
        mult_lsb_n125) );
  XOR2_X1 mult_lsb_U93 ( .A(mult_lsb_n40), .B(mult_lsb_n39), .Z(mult_lsb_n126)
         );
  XNOR2_X1 mult_lsb_U92 ( .A(mult_lsb_n124), .B(mult_lsb_n123), .ZN(
        InvUnmappedxD[25]) );
  XNOR2_X1 mult_lsb_U91 ( .A(mult_lsb_n42), .B(mult_lsb_n41), .ZN(
        mult_lsb_n123) );
  XOR2_X1 mult_lsb_U90 ( .A(mult_lsb_n44), .B(mult_lsb_n43), .Z(mult_lsb_n124)
         );
  XNOR2_X1 mult_lsb_U89 ( .A(mult_lsb_n122), .B(mult_lsb_n121), .ZN(
        InvUnmappedxD[24]) );
  XNOR2_X1 mult_lsb_U88 ( .A(mult_lsb_n46), .B(mult_lsb_n45), .ZN(
        mult_lsb_n121) );
  XOR2_X1 mult_lsb_U87 ( .A(mult_lsb_n48), .B(mult_lsb_n47), .Z(mult_lsb_n122)
         );
  XNOR2_X1 mult_lsb_U86 ( .A(mult_lsb_n120), .B(mult_lsb_n119), .ZN(
        InvUnmappedxD[19]) );
  XNOR2_X1 mult_lsb_U85 ( .A(mult_lsb_n50), .B(mult_lsb_n49), .ZN(
        mult_lsb_n119) );
  XOR2_X1 mult_lsb_U84 ( .A(mult_lsb_n52), .B(mult_lsb_n51), .Z(mult_lsb_n120)
         );
  XNOR2_X1 mult_lsb_U83 ( .A(mult_lsb_n118), .B(mult_lsb_n117), .ZN(
        InvUnmappedxD[18]) );
  XNOR2_X1 mult_lsb_U82 ( .A(mult_lsb_n54), .B(mult_lsb_n53), .ZN(
        mult_lsb_n117) );
  XOR2_X1 mult_lsb_U81 ( .A(mult_lsb_n56), .B(mult_lsb_n55), .Z(mult_lsb_n118)
         );
  XNOR2_X1 mult_lsb_U80 ( .A(mult_lsb_n116), .B(mult_lsb_n115), .ZN(
        InvUnmappedxD[17]) );
  XNOR2_X1 mult_lsb_U79 ( .A(mult_lsb_n58), .B(mult_lsb_n57), .ZN(
        mult_lsb_n115) );
  XOR2_X1 mult_lsb_U78 ( .A(mult_lsb_n60), .B(mult_lsb_n59), .Z(mult_lsb_n116)
         );
  XNOR2_X1 mult_lsb_U77 ( .A(mult_lsb_n114), .B(mult_lsb_n113), .ZN(
        InvUnmappedxD[16]) );
  XNOR2_X1 mult_lsb_U76 ( .A(mult_lsb_n62), .B(mult_lsb_n61), .ZN(
        mult_lsb_n113) );
  XOR2_X1 mult_lsb_U75 ( .A(mult_lsb_n64), .B(mult_lsb_n63), .Z(mult_lsb_n114)
         );
  XNOR2_X1 mult_lsb_U74 ( .A(mult_lsb_n112), .B(mult_lsb_n111), .ZN(
        InvUnmappedxD[11]) );
  XNOR2_X1 mult_lsb_U73 ( .A(mult_lsb_n66), .B(mult_lsb_n65), .ZN(
        mult_lsb_n111) );
  XOR2_X1 mult_lsb_U72 ( .A(mult_lsb_n68), .B(mult_lsb_n67), .Z(mult_lsb_n112)
         );
  XNOR2_X1 mult_lsb_U71 ( .A(mult_lsb_n110), .B(mult_lsb_n109), .ZN(
        InvUnmappedxD[10]) );
  XNOR2_X1 mult_lsb_U70 ( .A(mult_lsb_n70), .B(mult_lsb_n69), .ZN(
        mult_lsb_n109) );
  XOR2_X1 mult_lsb_U69 ( .A(mult_lsb_n72), .B(mult_lsb_n71), .Z(mult_lsb_n110)
         );
  XNOR2_X1 mult_lsb_U68 ( .A(mult_lsb_n108), .B(mult_lsb_n107), .ZN(
        InvUnmappedxD[9]) );
  XNOR2_X1 mult_lsb_U67 ( .A(mult_lsb_n74), .B(mult_lsb_n73), .ZN(
        mult_lsb_n107) );
  XOR2_X1 mult_lsb_U66 ( .A(mult_lsb_n76), .B(mult_lsb_n75), .Z(mult_lsb_n108)
         );
  XNOR2_X1 mult_lsb_U65 ( .A(mult_lsb_n106), .B(mult_lsb_n105), .ZN(
        InvUnmappedxD[8]) );
  XNOR2_X1 mult_lsb_U64 ( .A(mult_lsb_n78), .B(mult_lsb_n77), .ZN(
        mult_lsb_n105) );
  XOR2_X1 mult_lsb_U63 ( .A(mult_lsb_n80), .B(mult_lsb_n79), .Z(mult_lsb_n106)
         );
  XNOR2_X1 mult_lsb_U62 ( .A(mult_lsb_n104), .B(mult_lsb_n103), .ZN(
        InvUnmappedxD[3]) );
  XNOR2_X1 mult_lsb_U61 ( .A(mult_lsb_n82), .B(mult_lsb_n81), .ZN(
        mult_lsb_n103) );
  XOR2_X1 mult_lsb_U60 ( .A(mult_lsb_n84), .B(mult_lsb_n83), .Z(mult_lsb_n104)
         );
  XNOR2_X1 mult_lsb_U59 ( .A(mult_lsb_n102), .B(mult_lsb_n101), .ZN(
        InvUnmappedxD[2]) );
  XNOR2_X1 mult_lsb_U58 ( .A(mult_lsb_n86), .B(mult_lsb_n85), .ZN(
        mult_lsb_n101) );
  XOR2_X1 mult_lsb_U57 ( .A(mult_lsb_n88), .B(mult_lsb_n87), .Z(mult_lsb_n102)
         );
  XNOR2_X1 mult_lsb_U56 ( .A(mult_lsb_n100), .B(mult_lsb_n99), .ZN(
        InvUnmappedxD[1]) );
  XNOR2_X1 mult_lsb_U55 ( .A(mult_lsb_n90), .B(mult_lsb_n89), .ZN(mult_lsb_n99) );
  XOR2_X1 mult_lsb_U54 ( .A(mult_lsb_n92), .B(mult_lsb_n91), .Z(mult_lsb_n100)
         );
  XNOR2_X1 mult_lsb_U53 ( .A(mult_lsb_n98), .B(mult_lsb_n97), .ZN(
        InvUnmappedxD[0]) );
  XNOR2_X1 mult_lsb_U52 ( .A(mult_lsb_n94), .B(mult_lsb_n93), .ZN(mult_lsb_n97) );
  XOR2_X1 mult_lsb_U51 ( .A(mult_lsb_n96), .B(mult_lsb_n95), .Z(mult_lsb_n98)
         );
  XOR2_X1 mult_lsb_U50 ( .A(Zmul3xDI[11]), .B(mult_lsb_Xi_mul_Yj_9__3_), .Z(
        mult_lsb_FFxDN[39]) );
  XOR2_X1 mult_lsb_U49 ( .A(Zmul3xDI[10]), .B(mult_lsb_Xi_mul_Yj_9__2_), .Z(
        mult_lsb_FFxDN[38]) );
  XOR2_X1 mult_lsb_U48 ( .A(Zmul3xDI[9]), .B(mult_lsb_Xi_mul_Yj_9__1_), .Z(
        mult_lsb_FFxDN[37]) );
  XOR2_X1 mult_lsb_U47 ( .A(Zmul3xDI[8]), .B(mult_lsb_Xi_mul_Yj_9__0_), .Z(
        mult_lsb_FFxDN[36]) );
  XOR2_X1 mult_lsb_U46 ( .A(Zmul3xDI[7]), .B(mult_lsb_Xi_mul_Yj_8__3_), .Z(
        mult_lsb_FFxDN[35]) );
  XOR2_X1 mult_lsb_U45 ( .A(Zmul3xDI[6]), .B(mult_lsb_Xi_mul_Yj_8__2_), .Z(
        mult_lsb_FFxDN[34]) );
  XOR2_X1 mult_lsb_U44 ( .A(Zmul3xDI[5]), .B(mult_lsb_Xi_mul_Yj_8__1_), .Z(
        mult_lsb_FFxDN[33]) );
  XOR2_X1 mult_lsb_U43 ( .A(Zmul3xDI[4]), .B(mult_lsb_Xi_mul_Yj_8__0_), .Z(
        mult_lsb_FFxDN[32]) );
  XOR2_X1 mult_lsb_U42 ( .A(Zmul3xDI[19]), .B(mult_lsb_Xi_mul_Yj_7__3_), .Z(
        mult_lsb_FFxDN[31]) );
  XOR2_X1 mult_lsb_U41 ( .A(Zmul3xDI[18]), .B(mult_lsb_Xi_mul_Yj_7__2_), .Z(
        mult_lsb_FFxDN[30]) );
  XOR2_X1 mult_lsb_U40 ( .A(Zmul3xDI[17]), .B(mult_lsb_Xi_mul_Yj_7__1_), .Z(
        mult_lsb_FFxDN[29]) );
  XOR2_X1 mult_lsb_U39 ( .A(Zmul3xDI[16]), .B(mult_lsb_Xi_mul_Yj_7__0_), .Z(
        mult_lsb_FFxDN[28]) );
  XOR2_X1 mult_lsb_U38 ( .A(Zmul3xDI[11]), .B(mult_lsb_Xi_mul_Yj_6__3_), .Z(
        mult_lsb_FFxDN[27]) );
  XOR2_X1 mult_lsb_U37 ( .A(Zmul3xDI[10]), .B(mult_lsb_Xi_mul_Yj_6__2_), .Z(
        mult_lsb_FFxDN[26]) );
  XOR2_X1 mult_lsb_U36 ( .A(Zmul3xDI[9]), .B(mult_lsb_Xi_mul_Yj_6__1_), .Z(
        mult_lsb_FFxDN[25]) );
  XOR2_X1 mult_lsb_U35 ( .A(Zmul3xDI[8]), .B(mult_lsb_Xi_mul_Yj_6__0_), .Z(
        mult_lsb_FFxDN[24]) );
  XOR2_X1 mult_lsb_U34 ( .A(Zmul3xDI[3]), .B(mult_lsb_Xi_mul_Yj_4__3_), .Z(
        mult_lsb_FFxDN[19]) );
  XOR2_X1 mult_lsb_U33 ( .A(Zmul3xDI[2]), .B(mult_lsb_Xi_mul_Yj_4__2_), .Z(
        mult_lsb_FFxDN[18]) );
  XOR2_X1 mult_lsb_U32 ( .A(Zmul3xDI[1]), .B(mult_lsb_Xi_mul_Yj_4__1_), .Z(
        mult_lsb_FFxDN[17]) );
  XOR2_X1 mult_lsb_U31 ( .A(Zmul3xDI[0]), .B(mult_lsb_Xi_mul_Yj_4__0_), .Z(
        mult_lsb_FFxDN[16]) );
  XOR2_X1 mult_lsb_U30 ( .A(Zmul3xDI[15]), .B(mult_lsb_Xi_mul_Yj_3__3_), .Z(
        mult_lsb_FFxDN[15]) );
  XOR2_X1 mult_lsb_U29 ( .A(Zmul3xDI[14]), .B(mult_lsb_Xi_mul_Yj_3__2_), .Z(
        mult_lsb_FFxDN[14]) );
  XOR2_X1 mult_lsb_U28 ( .A(Zmul3xDI[13]), .B(mult_lsb_Xi_mul_Yj_3__1_), .Z(
        mult_lsb_FFxDN[13]) );
  XOR2_X1 mult_lsb_U27 ( .A(Zmul3xDI[12]), .B(mult_lsb_Xi_mul_Yj_3__0_), .Z(
        mult_lsb_FFxDN[12]) );
  XOR2_X1 mult_lsb_U26 ( .A(Zmul3xDI[7]), .B(mult_lsb_Xi_mul_Yj_2__3_), .Z(
        mult_lsb_FFxDN[11]) );
  XOR2_X1 mult_lsb_U25 ( .A(Zmul3xDI[6]), .B(mult_lsb_Xi_mul_Yj_2__2_), .Z(
        mult_lsb_FFxDN[10]) );
  XOR2_X1 mult_lsb_U24 ( .A(Zmul3xDI[5]), .B(mult_lsb_Xi_mul_Yj_2__1_), .Z(
        mult_lsb_FFxDN[9]) );
  XOR2_X1 mult_lsb_U23 ( .A(Zmul3xDI[4]), .B(mult_lsb_Xi_mul_Yj_2__0_), .Z(
        mult_lsb_FFxDN[8]) );
  XOR2_X1 mult_lsb_U22 ( .A(Zmul3xDI[3]), .B(mult_lsb_Xi_mul_Yj_1__3_), .Z(
        mult_lsb_FFxDN[7]) );
  XOR2_X1 mult_lsb_U21 ( .A(Zmul3xDI[2]), .B(mult_lsb_Xi_mul_Yj_1__2_), .Z(
        mult_lsb_FFxDN[6]) );
  XOR2_X1 mult_lsb_U20 ( .A(Zmul3xDI[1]), .B(mult_lsb_Xi_mul_Yj_1__1_), .Z(
        mult_lsb_FFxDN[5]) );
  XOR2_X1 mult_lsb_U19 ( .A(Zmul3xDI[0]), .B(mult_lsb_Xi_mul_Yj_1__0_), .Z(
        mult_lsb_FFxDN[4]) );
  XOR2_X1 mult_lsb_U18 ( .A(Zmul3xDI[23]), .B(mult_lsb_Xi_mul_Yj_14__3_), .Z(
        mult_lsb_FFxDN[59]) );
  XOR2_X1 mult_lsb_U17 ( .A(Zmul3xDI[22]), .B(mult_lsb_Xi_mul_Yj_14__2_), .Z(
        mult_lsb_FFxDN[58]) );
  XOR2_X1 mult_lsb_U16 ( .A(Zmul3xDI[21]), .B(mult_lsb_Xi_mul_Yj_14__1_), .Z(
        mult_lsb_FFxDN[57]) );
  XOR2_X1 mult_lsb_U15 ( .A(Zmul3xDI[20]), .B(mult_lsb_Xi_mul_Yj_14__0_), .Z(
        mult_lsb_FFxDN[56]) );
  XOR2_X1 mult_lsb_U14 ( .A(Zmul3xDI[19]), .B(mult_lsb_Xi_mul_Yj_13__3_), .Z(
        mult_lsb_FFxDN[55]) );
  XOR2_X1 mult_lsb_U13 ( .A(Zmul3xDI[18]), .B(mult_lsb_Xi_mul_Yj_13__2_), .Z(
        mult_lsb_FFxDN[54]) );
  XOR2_X1 mult_lsb_U12 ( .A(Zmul3xDI[17]), .B(mult_lsb_Xi_mul_Yj_13__1_), .Z(
        mult_lsb_FFxDN[53]) );
  XOR2_X1 mult_lsb_U11 ( .A(Zmul3xDI[16]), .B(mult_lsb_Xi_mul_Yj_13__0_), .Z(
        mult_lsb_FFxDN[52]) );
  XOR2_X1 mult_lsb_U10 ( .A(Zmul3xDI[15]), .B(mult_lsb_Xi_mul_Yj_12__3_), .Z(
        mult_lsb_FFxDN[51]) );
  XOR2_X1 mult_lsb_U9 ( .A(Zmul3xDI[14]), .B(mult_lsb_Xi_mul_Yj_12__2_), .Z(
        mult_lsb_FFxDN[50]) );
  XOR2_X1 mult_lsb_U8 ( .A(Zmul3xDI[13]), .B(mult_lsb_Xi_mul_Yj_12__1_), .Z(
        mult_lsb_FFxDN[49]) );
  XOR2_X1 mult_lsb_U7 ( .A(Zmul3xDI[12]), .B(mult_lsb_Xi_mul_Yj_12__0_), .Z(
        mult_lsb_FFxDN[48]) );
  XOR2_X1 mult_lsb_U6 ( .A(Zmul3xDI[23]), .B(mult_lsb_Xi_mul_Yj_11__3_), .Z(
        mult_lsb_FFxDN[47]) );
  XOR2_X1 mult_lsb_U5 ( .A(Zmul3xDI[22]), .B(mult_lsb_Xi_mul_Yj_11__2_), .Z(
        mult_lsb_FFxDN[46]) );
  XOR2_X1 mult_lsb_U4 ( .A(Zmul3xDI[21]), .B(mult_lsb_Xi_mul_Yj_11__1_), .Z(
        mult_lsb_FFxDN[45]) );
  XOR2_X1 mult_lsb_U3 ( .A(Zmul3xDI[20]), .B(mult_lsb_Xi_mul_Yj_11__0_), .Z(
        mult_lsb_FFxDN[44]) );
  DFF_X1 mult_lsb_FFxDP_reg_1__3_ ( .D(mult_lsb_FFxDN[7]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n84) );
  DFF_X1 mult_lsb_FFxDP_reg_2__3_ ( .D(mult_lsb_FFxDN[11]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n81) );
  DFF_X1 mult_lsb_FFxDP_reg_3__3_ ( .D(mult_lsb_FFxDN[15]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n82) );
  DFF_X1 mult_lsb_FFxDP_reg_4__3_ ( .D(mult_lsb_FFxDN[19]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n67) );
  DFF_X1 mult_lsb_FFxDP_reg_6__3_ ( .D(mult_lsb_FFxDN[27]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n65) );
  DFF_X1 mult_lsb_FFxDP_reg_7__3_ ( .D(mult_lsb_FFxDN[31]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n66) );
  DFF_X1 mult_lsb_FFxDP_reg_8__3_ ( .D(mult_lsb_FFxDN[35]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n49) );
  DFF_X1 mult_lsb_FFxDP_reg_9__3_ ( .D(mult_lsb_FFxDN[39]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n50) );
  DFF_X1 mult_lsb_FFxDP_reg_11__3_ ( .D(mult_lsb_FFxDN[47]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n52) );
  DFF_X1 mult_lsb_FFxDP_reg_12__3_ ( .D(mult_lsb_FFxDN[51]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n35) );
  DFF_X1 mult_lsb_FFxDP_reg_13__3_ ( .D(mult_lsb_FFxDN[55]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n36) );
  DFF_X1 mult_lsb_FFxDP_reg_14__3_ ( .D(mult_lsb_FFxDN[59]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n33) );
  DFF_X1 mult_lsb_FFxDP_reg_1__1_ ( .D(mult_lsb_FFxDN[5]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n92) );
  DFF_X1 mult_lsb_FFxDP_reg_2__1_ ( .D(mult_lsb_FFxDN[9]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n89) );
  DFF_X1 mult_lsb_FFxDP_reg_3__1_ ( .D(mult_lsb_FFxDN[13]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n90) );
  DFF_X1 mult_lsb_FFxDP_reg_4__1_ ( .D(mult_lsb_FFxDN[17]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n75) );
  DFF_X1 mult_lsb_FFxDP_reg_6__1_ ( .D(mult_lsb_FFxDN[25]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n73) );
  DFF_X1 mult_lsb_FFxDP_reg_7__1_ ( .D(mult_lsb_FFxDN[29]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n74) );
  DFF_X1 mult_lsb_FFxDP_reg_8__1_ ( .D(mult_lsb_FFxDN[33]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n57) );
  DFF_X1 mult_lsb_FFxDP_reg_9__1_ ( .D(mult_lsb_FFxDN[37]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n58) );
  DFF_X1 mult_lsb_FFxDP_reg_11__1_ ( .D(mult_lsb_FFxDN[45]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n60) );
  DFF_X1 mult_lsb_FFxDP_reg_12__1_ ( .D(mult_lsb_FFxDN[49]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n43) );
  DFF_X1 mult_lsb_FFxDP_reg_13__1_ ( .D(mult_lsb_FFxDN[53]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n44) );
  DFF_X1 mult_lsb_FFxDP_reg_14__1_ ( .D(mult_lsb_FFxDN[57]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n41) );
  DFF_X1 mult_lsb_FFxDP_reg_1__2_ ( .D(mult_lsb_FFxDN[6]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n88) );
  DFF_X1 mult_lsb_FFxDP_reg_2__2_ ( .D(mult_lsb_FFxDN[10]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n85) );
  DFF_X1 mult_lsb_FFxDP_reg_3__2_ ( .D(mult_lsb_FFxDN[14]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n86) );
  DFF_X1 mult_lsb_FFxDP_reg_4__2_ ( .D(mult_lsb_FFxDN[18]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n71) );
  DFF_X1 mult_lsb_FFxDP_reg_6__2_ ( .D(mult_lsb_FFxDN[26]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n69) );
  DFF_X1 mult_lsb_FFxDP_reg_7__2_ ( .D(mult_lsb_FFxDN[30]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n70) );
  DFF_X1 mult_lsb_FFxDP_reg_8__2_ ( .D(mult_lsb_FFxDN[34]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n53) );
  DFF_X1 mult_lsb_FFxDP_reg_9__2_ ( .D(mult_lsb_FFxDN[38]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n54) );
  DFF_X1 mult_lsb_FFxDP_reg_11__2_ ( .D(mult_lsb_FFxDN[46]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n56) );
  DFF_X1 mult_lsb_FFxDP_reg_12__2_ ( .D(mult_lsb_FFxDN[50]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n39) );
  DFF_X1 mult_lsb_FFxDP_reg_13__2_ ( .D(mult_lsb_FFxDN[54]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n40) );
  DFF_X1 mult_lsb_FFxDP_reg_14__2_ ( .D(mult_lsb_FFxDN[58]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n37) );
  DFF_X1 mult_lsb_FFxDP_reg_1__0_ ( .D(mult_lsb_FFxDN[4]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n96) );
  DFF_X1 mult_lsb_FFxDP_reg_2__0_ ( .D(mult_lsb_FFxDN[8]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n93) );
  DFF_X1 mult_lsb_FFxDP_reg_3__0_ ( .D(mult_lsb_FFxDN[12]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n94) );
  DFF_X1 mult_lsb_FFxDP_reg_4__0_ ( .D(mult_lsb_FFxDN[16]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n79) );
  DFF_X1 mult_lsb_FFxDP_reg_6__0_ ( .D(mult_lsb_FFxDN[24]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n77) );
  DFF_X1 mult_lsb_FFxDP_reg_7__0_ ( .D(mult_lsb_FFxDN[28]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n78) );
  DFF_X1 mult_lsb_FFxDP_reg_8__0_ ( .D(mult_lsb_FFxDN[32]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n61) );
  DFF_X1 mult_lsb_FFxDP_reg_9__0_ ( .D(mult_lsb_FFxDN[36]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n62) );
  DFF_X1 mult_lsb_FFxDP_reg_11__0_ ( .D(mult_lsb_FFxDN[44]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n64) );
  DFF_X1 mult_lsb_FFxDP_reg_12__0_ ( .D(mult_lsb_FFxDN[48]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n47) );
  DFF_X1 mult_lsb_FFxDP_reg_13__0_ ( .D(mult_lsb_FFxDN[52]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n48) );
  DFF_X1 mult_lsb_FFxDP_reg_14__0_ ( .D(mult_lsb_FFxDN[56]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n45) );
  DFF_X1 mult_lsb_FFxDP_reg_0__3_ ( .D(mult_lsb_FFxDN[3]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n83) );
  DFF_X1 mult_lsb_FFxDP_reg_5__3_ ( .D(mult_lsb_FFxDN[23]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n68) );
  DFF_X1 mult_lsb_FFxDP_reg_10__3_ ( .D(mult_lsb_FFxDN[43]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n51) );
  DFF_X1 mult_lsb_FFxDP_reg_15__3_ ( .D(mult_lsb_FFxDN[63]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n34) );
  DFF_X1 mult_lsb_FFxDP_reg_0__1_ ( .D(mult_lsb_FFxDN[1]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n91) );
  DFF_X1 mult_lsb_FFxDP_reg_5__1_ ( .D(mult_lsb_FFxDN[21]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n76) );
  DFF_X1 mult_lsb_FFxDP_reg_10__1_ ( .D(mult_lsb_FFxDN[41]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n59) );
  DFF_X1 mult_lsb_FFxDP_reg_15__1_ ( .D(mult_lsb_FFxDN[61]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n42) );
  DFF_X1 mult_lsb_FFxDP_reg_0__2_ ( .D(mult_lsb_FFxDN[2]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n87) );
  DFF_X1 mult_lsb_FFxDP_reg_5__2_ ( .D(mult_lsb_FFxDN[22]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n72) );
  DFF_X1 mult_lsb_FFxDP_reg_10__2_ ( .D(mult_lsb_FFxDN[42]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n55) );
  DFF_X1 mult_lsb_FFxDP_reg_15__2_ ( .D(mult_lsb_FFxDN[62]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n38) );
  DFF_X1 mult_lsb_FFxDP_reg_0__0_ ( .D(mult_lsb_FFxDN[0]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n95) );
  DFF_X1 mult_lsb_FFxDP_reg_5__0_ ( .D(mult_lsb_FFxDN[20]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n80) );
  DFF_X1 mult_lsb_FFxDP_reg_10__0_ ( .D(mult_lsb_FFxDN[40]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n63) );
  DFF_X1 mult_lsb_FFxDP_reg_15__0_ ( .D(mult_lsb_FFxDN[60]), .CK(ClkxCI), .Q(), 
        .QN(mult_lsb_n46) );
  XNOR2_X1 mult_lsb_gf4_mul_3_3_U29 ( .A(mult_lsb_gf4_mul_3_3_n77), .B(
        mult_lsb_gf4_mul_3_3_n76), .ZN(mult_lsb_FFxDN[63]) );
  NAND2_X1 mult_lsb_gf4_mul_3_3_U28 ( .A1(n119), .A2(Y1_4xDP[15]), .ZN(
        mult_lsb_gf4_mul_3_3_n76) );
  XOR2_X1 mult_lsb_gf4_mul_3_3_U27 ( .A(mult_lsb_gf4_mul_3_3_n75), .B(
        mult_lsb_gf4_mul_3_3_n74), .Z(mult_lsb_gf4_mul_3_3_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_3_3_U26 ( .A(mult_lsb_gf4_mul_3_3_n73), .B(
        mult_lsb_gf4_mul_3_3_n72), .ZN(mult_lsb_FFxDN[62]) );
  NAND2_X1 mult_lsb_gf4_mul_3_3_U25 ( .A1(n117), .A2(Y1_4xDP[14]), .ZN(
        mult_lsb_gf4_mul_3_3_n72) );
  XOR2_X1 mult_lsb_gf4_mul_3_3_U24 ( .A(mult_lsb_gf4_mul_3_3_n74), .B(
        mult_lsb_gf4_mul_3_3_n71), .Z(mult_lsb_gf4_mul_3_3_n73) );
  NOR2_X1 mult_lsb_gf4_mul_3_3_U23 ( .A1(mult_lsb_gf4_mul_3_3_n70), .A2(
        mult_lsb_gf4_mul_3_3_n69), .ZN(mult_lsb_gf4_mul_3_3_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_3_3_U22 ( .A(n117), .B(n119), .ZN(
        mult_lsb_gf4_mul_3_3_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_3_3_U21 ( .A(Y1_4xDP[14]), .B(Y1_4xDP[15]), .ZN(
        mult_lsb_gf4_mul_3_3_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_3_3_U20 ( .A(mult_lsb_gf4_mul_3_3_n68), .B(
        mult_lsb_gf4_mul_3_3_n67), .ZN(mult_lsb_FFxDN[61]) );
  NAND2_X1 mult_lsb_gf4_mul_3_3_U19 ( .A1(n115), .A2(Y1_4xDP[13]), .ZN(
        mult_lsb_gf4_mul_3_3_n67) );
  XOR2_X1 mult_lsb_gf4_mul_3_3_U18 ( .A(mult_lsb_gf4_mul_3_3_n75), .B(
        mult_lsb_gf4_mul_3_3_n66), .Z(mult_lsb_gf4_mul_3_3_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_3_3_U17 ( .A(mult_lsb_gf4_mul_3_3_n65), .B(
        mult_lsb_gf4_mul_3_3_n64), .ZN(mult_lsb_gf4_mul_3_3_n75) );
  NAND2_X1 mult_lsb_gf4_mul_3_3_U16 ( .A1(mult_lsb_gf4_mul_3_3_n63), .A2(
        mult_lsb_gf4_mul_3_3_n62), .ZN(mult_lsb_gf4_mul_3_3_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_3_3_U15 ( .A(mult_lsb_gf4_mul_3_3_n61), .B(
        mult_lsb_gf4_mul_3_3_n60), .ZN(mult_lsb_gf4_mul_3_3_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_3_3_U14 ( .A(mult_lsb_gf4_mul_3_3_n59), .B(
        mult_lsb_gf4_mul_3_3_n58), .ZN(mult_lsb_gf4_mul_3_3_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_3_3_U13 ( .A(mult_lsb_gf4_mul_3_3_n57), .B(
        mult_lsb_gf4_mul_3_3_n56), .ZN(mult_lsb_FFxDN[60]) );
  NAND2_X1 mult_lsb_gf4_mul_3_3_U12 ( .A1(n113), .A2(Y1_4xDP[12]), .ZN(
        mult_lsb_gf4_mul_3_3_n56) );
  XOR2_X1 mult_lsb_gf4_mul_3_3_U11 ( .A(mult_lsb_gf4_mul_3_3_n66), .B(
        mult_lsb_gf4_mul_3_3_n71), .Z(mult_lsb_gf4_mul_3_3_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_3_3_U10 ( .A(mult_lsb_gf4_mul_3_3_n55), .B(
        mult_lsb_gf4_mul_3_3_n65), .ZN(mult_lsb_gf4_mul_3_3_n71) );
  NOR2_X1 mult_lsb_gf4_mul_3_3_U9 ( .A1(mult_lsb_gf4_mul_3_3_n61), .A2(
        mult_lsb_gf4_mul_3_3_n59), .ZN(mult_lsb_gf4_mul_3_3_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_3_3_U8 ( .A(n113), .B(n117), .ZN(
        mult_lsb_gf4_mul_3_3_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_3_3_U7 ( .A(Y1_4xDP[12]), .B(Y1_4xDP[14]), .ZN(
        mult_lsb_gf4_mul_3_3_n61) );
  NAND2_X1 mult_lsb_gf4_mul_3_3_U6 ( .A1(mult_lsb_gf4_mul_3_3_n58), .A2(
        mult_lsb_gf4_mul_3_3_n60), .ZN(mult_lsb_gf4_mul_3_3_n55) );
  XOR2_X1 mult_lsb_gf4_mul_3_3_U5 ( .A(Y1_4xDP[13]), .B(Y1_4xDP[15]), .Z(
        mult_lsb_gf4_mul_3_3_n60) );
  XOR2_X1 mult_lsb_gf4_mul_3_3_U4 ( .A(n115), .B(n119), .Z(
        mult_lsb_gf4_mul_3_3_n58) );
  NOR2_X1 mult_lsb_gf4_mul_3_3_U3 ( .A1(mult_lsb_gf4_mul_3_3_n54), .A2(
        mult_lsb_gf4_mul_3_3_n53), .ZN(mult_lsb_gf4_mul_3_3_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_3_3_U2 ( .A(n113), .B(n115), .ZN(
        mult_lsb_gf4_mul_3_3_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_3_3_U1 ( .A(Y1_4xDP[12]), .B(Y1_4xDP[13]), .ZN(
        mult_lsb_gf4_mul_3_3_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_3_2_U29 ( .A(mult_lsb_gf4_mul_3_2_n77), .B(
        mult_lsb_gf4_mul_3_2_n76), .ZN(mult_lsb_Xi_mul_Yj_14__3_) );
  NAND2_X1 mult_lsb_gf4_mul_3_2_U28 ( .A1(n119), .A2(Y1_4xDP[11]), .ZN(
        mult_lsb_gf4_mul_3_2_n76) );
  XOR2_X1 mult_lsb_gf4_mul_3_2_U27 ( .A(mult_lsb_gf4_mul_3_2_n75), .B(
        mult_lsb_gf4_mul_3_2_n74), .Z(mult_lsb_gf4_mul_3_2_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_3_2_U26 ( .A(mult_lsb_gf4_mul_3_2_n73), .B(
        mult_lsb_gf4_mul_3_2_n72), .ZN(mult_lsb_Xi_mul_Yj_14__2_) );
  NAND2_X1 mult_lsb_gf4_mul_3_2_U25 ( .A1(n117), .A2(Y1_4xDP[10]), .ZN(
        mult_lsb_gf4_mul_3_2_n72) );
  XOR2_X1 mult_lsb_gf4_mul_3_2_U24 ( .A(mult_lsb_gf4_mul_3_2_n74), .B(
        mult_lsb_gf4_mul_3_2_n71), .Z(mult_lsb_gf4_mul_3_2_n73) );
  NOR2_X1 mult_lsb_gf4_mul_3_2_U23 ( .A1(mult_lsb_gf4_mul_3_2_n70), .A2(
        mult_lsb_gf4_mul_3_2_n69), .ZN(mult_lsb_gf4_mul_3_2_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_3_2_U22 ( .A(n117), .B(n119), .ZN(
        mult_lsb_gf4_mul_3_2_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_3_2_U21 ( .A(Y1_4xDP[10]), .B(Y1_4xDP[11]), .ZN(
        mult_lsb_gf4_mul_3_2_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_3_2_U20 ( .A(mult_lsb_gf4_mul_3_2_n68), .B(
        mult_lsb_gf4_mul_3_2_n67), .ZN(mult_lsb_Xi_mul_Yj_14__1_) );
  NAND2_X1 mult_lsb_gf4_mul_3_2_U19 ( .A1(n115), .A2(Y1_4xDP[9]), .ZN(
        mult_lsb_gf4_mul_3_2_n67) );
  XOR2_X1 mult_lsb_gf4_mul_3_2_U18 ( .A(mult_lsb_gf4_mul_3_2_n75), .B(
        mult_lsb_gf4_mul_3_2_n66), .Z(mult_lsb_gf4_mul_3_2_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_3_2_U17 ( .A(mult_lsb_gf4_mul_3_2_n65), .B(
        mult_lsb_gf4_mul_3_2_n64), .ZN(mult_lsb_gf4_mul_3_2_n75) );
  NAND2_X1 mult_lsb_gf4_mul_3_2_U16 ( .A1(mult_lsb_gf4_mul_3_2_n63), .A2(
        mult_lsb_gf4_mul_3_2_n62), .ZN(mult_lsb_gf4_mul_3_2_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_3_2_U15 ( .A(mult_lsb_gf4_mul_3_2_n61), .B(
        mult_lsb_gf4_mul_3_2_n60), .ZN(mult_lsb_gf4_mul_3_2_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_3_2_U14 ( .A(mult_lsb_gf4_mul_3_2_n59), .B(
        mult_lsb_gf4_mul_3_2_n58), .ZN(mult_lsb_gf4_mul_3_2_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_3_2_U13 ( .A(mult_lsb_gf4_mul_3_2_n57), .B(
        mult_lsb_gf4_mul_3_2_n56), .ZN(mult_lsb_Xi_mul_Yj_14__0_) );
  NAND2_X1 mult_lsb_gf4_mul_3_2_U12 ( .A1(n113), .A2(Y1_4xDP[8]), .ZN(
        mult_lsb_gf4_mul_3_2_n56) );
  XOR2_X1 mult_lsb_gf4_mul_3_2_U11 ( .A(mult_lsb_gf4_mul_3_2_n66), .B(
        mult_lsb_gf4_mul_3_2_n71), .Z(mult_lsb_gf4_mul_3_2_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_3_2_U10 ( .A(mult_lsb_gf4_mul_3_2_n55), .B(
        mult_lsb_gf4_mul_3_2_n65), .ZN(mult_lsb_gf4_mul_3_2_n71) );
  NOR2_X1 mult_lsb_gf4_mul_3_2_U9 ( .A1(mult_lsb_gf4_mul_3_2_n61), .A2(
        mult_lsb_gf4_mul_3_2_n59), .ZN(mult_lsb_gf4_mul_3_2_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_3_2_U8 ( .A(n113), .B(n117), .ZN(
        mult_lsb_gf4_mul_3_2_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_3_2_U7 ( .A(Y1_4xDP[8]), .B(Y1_4xDP[10]), .ZN(
        mult_lsb_gf4_mul_3_2_n61) );
  NAND2_X1 mult_lsb_gf4_mul_3_2_U6 ( .A1(mult_lsb_gf4_mul_3_2_n58), .A2(
        mult_lsb_gf4_mul_3_2_n60), .ZN(mult_lsb_gf4_mul_3_2_n55) );
  XOR2_X1 mult_lsb_gf4_mul_3_2_U5 ( .A(Y1_4xDP[9]), .B(Y1_4xDP[11]), .Z(
        mult_lsb_gf4_mul_3_2_n60) );
  XOR2_X1 mult_lsb_gf4_mul_3_2_U4 ( .A(n115), .B(n119), .Z(
        mult_lsb_gf4_mul_3_2_n58) );
  NOR2_X1 mult_lsb_gf4_mul_3_2_U3 ( .A1(mult_lsb_gf4_mul_3_2_n54), .A2(
        mult_lsb_gf4_mul_3_2_n53), .ZN(mult_lsb_gf4_mul_3_2_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_3_2_U2 ( .A(n113), .B(n115), .ZN(
        mult_lsb_gf4_mul_3_2_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_3_2_U1 ( .A(Y1_4xDP[8]), .B(Y1_4xDP[9]), .ZN(
        mult_lsb_gf4_mul_3_2_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_3_1_U29 ( .A(mult_lsb_gf4_mul_3_1_n77), .B(
        mult_lsb_gf4_mul_3_1_n76), .ZN(mult_lsb_Xi_mul_Yj_13__3_) );
  NAND2_X1 mult_lsb_gf4_mul_3_1_U28 ( .A1(n119), .A2(Y1_4xDP[7]), .ZN(
        mult_lsb_gf4_mul_3_1_n76) );
  XOR2_X1 mult_lsb_gf4_mul_3_1_U27 ( .A(mult_lsb_gf4_mul_3_1_n75), .B(
        mult_lsb_gf4_mul_3_1_n74), .Z(mult_lsb_gf4_mul_3_1_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_3_1_U26 ( .A(mult_lsb_gf4_mul_3_1_n73), .B(
        mult_lsb_gf4_mul_3_1_n72), .ZN(mult_lsb_Xi_mul_Yj_13__2_) );
  NAND2_X1 mult_lsb_gf4_mul_3_1_U25 ( .A1(n117), .A2(Y1_4xDP[6]), .ZN(
        mult_lsb_gf4_mul_3_1_n72) );
  XOR2_X1 mult_lsb_gf4_mul_3_1_U24 ( .A(mult_lsb_gf4_mul_3_1_n74), .B(
        mult_lsb_gf4_mul_3_1_n71), .Z(mult_lsb_gf4_mul_3_1_n73) );
  NOR2_X1 mult_lsb_gf4_mul_3_1_U23 ( .A1(mult_lsb_gf4_mul_3_1_n70), .A2(
        mult_lsb_gf4_mul_3_1_n69), .ZN(mult_lsb_gf4_mul_3_1_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_3_1_U22 ( .A(n117), .B(n119), .ZN(
        mult_lsb_gf4_mul_3_1_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_3_1_U21 ( .A(Y1_4xDP[6]), .B(Y1_4xDP[7]), .ZN(
        mult_lsb_gf4_mul_3_1_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_3_1_U20 ( .A(mult_lsb_gf4_mul_3_1_n68), .B(
        mult_lsb_gf4_mul_3_1_n67), .ZN(mult_lsb_Xi_mul_Yj_13__1_) );
  NAND2_X1 mult_lsb_gf4_mul_3_1_U19 ( .A1(n115), .A2(Y1_4xDP[5]), .ZN(
        mult_lsb_gf4_mul_3_1_n67) );
  XOR2_X1 mult_lsb_gf4_mul_3_1_U18 ( .A(mult_lsb_gf4_mul_3_1_n75), .B(
        mult_lsb_gf4_mul_3_1_n66), .Z(mult_lsb_gf4_mul_3_1_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_3_1_U17 ( .A(mult_lsb_gf4_mul_3_1_n65), .B(
        mult_lsb_gf4_mul_3_1_n64), .ZN(mult_lsb_gf4_mul_3_1_n75) );
  NAND2_X1 mult_lsb_gf4_mul_3_1_U16 ( .A1(mult_lsb_gf4_mul_3_1_n63), .A2(
        mult_lsb_gf4_mul_3_1_n62), .ZN(mult_lsb_gf4_mul_3_1_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_3_1_U15 ( .A(mult_lsb_gf4_mul_3_1_n61), .B(
        mult_lsb_gf4_mul_3_1_n60), .ZN(mult_lsb_gf4_mul_3_1_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_3_1_U14 ( .A(mult_lsb_gf4_mul_3_1_n59), .B(
        mult_lsb_gf4_mul_3_1_n58), .ZN(mult_lsb_gf4_mul_3_1_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_3_1_U13 ( .A(mult_lsb_gf4_mul_3_1_n57), .B(
        mult_lsb_gf4_mul_3_1_n56), .ZN(mult_lsb_Xi_mul_Yj_13__0_) );
  NAND2_X1 mult_lsb_gf4_mul_3_1_U12 ( .A1(n113), .A2(Y1_4xDP[4]), .ZN(
        mult_lsb_gf4_mul_3_1_n56) );
  XOR2_X1 mult_lsb_gf4_mul_3_1_U11 ( .A(mult_lsb_gf4_mul_3_1_n66), .B(
        mult_lsb_gf4_mul_3_1_n71), .Z(mult_lsb_gf4_mul_3_1_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_3_1_U10 ( .A(mult_lsb_gf4_mul_3_1_n55), .B(
        mult_lsb_gf4_mul_3_1_n65), .ZN(mult_lsb_gf4_mul_3_1_n71) );
  NOR2_X1 mult_lsb_gf4_mul_3_1_U9 ( .A1(mult_lsb_gf4_mul_3_1_n61), .A2(
        mult_lsb_gf4_mul_3_1_n59), .ZN(mult_lsb_gf4_mul_3_1_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_3_1_U8 ( .A(n113), .B(n117), .ZN(
        mult_lsb_gf4_mul_3_1_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_3_1_U7 ( .A(Y1_4xDP[4]), .B(Y1_4xDP[6]), .ZN(
        mult_lsb_gf4_mul_3_1_n61) );
  NAND2_X1 mult_lsb_gf4_mul_3_1_U6 ( .A1(mult_lsb_gf4_mul_3_1_n58), .A2(
        mult_lsb_gf4_mul_3_1_n60), .ZN(mult_lsb_gf4_mul_3_1_n55) );
  XOR2_X1 mult_lsb_gf4_mul_3_1_U5 ( .A(Y1_4xDP[5]), .B(Y1_4xDP[7]), .Z(
        mult_lsb_gf4_mul_3_1_n60) );
  XOR2_X1 mult_lsb_gf4_mul_3_1_U4 ( .A(n115), .B(n119), .Z(
        mult_lsb_gf4_mul_3_1_n58) );
  NOR2_X1 mult_lsb_gf4_mul_3_1_U3 ( .A1(mult_lsb_gf4_mul_3_1_n54), .A2(
        mult_lsb_gf4_mul_3_1_n53), .ZN(mult_lsb_gf4_mul_3_1_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_3_1_U2 ( .A(n113), .B(n115), .ZN(
        mult_lsb_gf4_mul_3_1_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_3_1_U1 ( .A(Y1_4xDP[4]), .B(Y1_4xDP[5]), .ZN(
        mult_lsb_gf4_mul_3_1_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_3_0_U29 ( .A(mult_lsb_gf4_mul_3_0_n77), .B(
        mult_lsb_gf4_mul_3_0_n76), .ZN(mult_lsb_Xi_mul_Yj_12__3_) );
  NAND2_X1 mult_lsb_gf4_mul_3_0_U28 ( .A1(n119), .A2(Y1_4xDP[3]), .ZN(
        mult_lsb_gf4_mul_3_0_n76) );
  XOR2_X1 mult_lsb_gf4_mul_3_0_U27 ( .A(mult_lsb_gf4_mul_3_0_n75), .B(
        mult_lsb_gf4_mul_3_0_n74), .Z(mult_lsb_gf4_mul_3_0_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_3_0_U26 ( .A(mult_lsb_gf4_mul_3_0_n73), .B(
        mult_lsb_gf4_mul_3_0_n72), .ZN(mult_lsb_Xi_mul_Yj_12__2_) );
  NAND2_X1 mult_lsb_gf4_mul_3_0_U25 ( .A1(n117), .A2(Y1_4xDP[2]), .ZN(
        mult_lsb_gf4_mul_3_0_n72) );
  XOR2_X1 mult_lsb_gf4_mul_3_0_U24 ( .A(mult_lsb_gf4_mul_3_0_n74), .B(
        mult_lsb_gf4_mul_3_0_n71), .Z(mult_lsb_gf4_mul_3_0_n73) );
  NOR2_X1 mult_lsb_gf4_mul_3_0_U23 ( .A1(mult_lsb_gf4_mul_3_0_n70), .A2(
        mult_lsb_gf4_mul_3_0_n69), .ZN(mult_lsb_gf4_mul_3_0_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_3_0_U22 ( .A(n117), .B(n119), .ZN(
        mult_lsb_gf4_mul_3_0_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_3_0_U21 ( .A(Y1_4xDP[2]), .B(Y1_4xDP[3]), .ZN(
        mult_lsb_gf4_mul_3_0_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_3_0_U20 ( .A(mult_lsb_gf4_mul_3_0_n68), .B(
        mult_lsb_gf4_mul_3_0_n67), .ZN(mult_lsb_Xi_mul_Yj_12__1_) );
  NAND2_X1 mult_lsb_gf4_mul_3_0_U19 ( .A1(n115), .A2(Y1_4xDP[1]), .ZN(
        mult_lsb_gf4_mul_3_0_n67) );
  XOR2_X1 mult_lsb_gf4_mul_3_0_U18 ( .A(mult_lsb_gf4_mul_3_0_n75), .B(
        mult_lsb_gf4_mul_3_0_n66), .Z(mult_lsb_gf4_mul_3_0_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_3_0_U17 ( .A(mult_lsb_gf4_mul_3_0_n65), .B(
        mult_lsb_gf4_mul_3_0_n64), .ZN(mult_lsb_gf4_mul_3_0_n75) );
  NAND2_X1 mult_lsb_gf4_mul_3_0_U16 ( .A1(mult_lsb_gf4_mul_3_0_n63), .A2(
        mult_lsb_gf4_mul_3_0_n62), .ZN(mult_lsb_gf4_mul_3_0_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_3_0_U15 ( .A(mult_lsb_gf4_mul_3_0_n61), .B(
        mult_lsb_gf4_mul_3_0_n60), .ZN(mult_lsb_gf4_mul_3_0_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_3_0_U14 ( .A(mult_lsb_gf4_mul_3_0_n59), .B(
        mult_lsb_gf4_mul_3_0_n58), .ZN(mult_lsb_gf4_mul_3_0_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_3_0_U13 ( .A(mult_lsb_gf4_mul_3_0_n57), .B(
        mult_lsb_gf4_mul_3_0_n56), .ZN(mult_lsb_Xi_mul_Yj_12__0_) );
  NAND2_X1 mult_lsb_gf4_mul_3_0_U12 ( .A1(n113), .A2(Y1_4xDP[0]), .ZN(
        mult_lsb_gf4_mul_3_0_n56) );
  XOR2_X1 mult_lsb_gf4_mul_3_0_U11 ( .A(mult_lsb_gf4_mul_3_0_n66), .B(
        mult_lsb_gf4_mul_3_0_n71), .Z(mult_lsb_gf4_mul_3_0_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_3_0_U10 ( .A(mult_lsb_gf4_mul_3_0_n55), .B(
        mult_lsb_gf4_mul_3_0_n65), .ZN(mult_lsb_gf4_mul_3_0_n71) );
  NOR2_X1 mult_lsb_gf4_mul_3_0_U9 ( .A1(mult_lsb_gf4_mul_3_0_n61), .A2(
        mult_lsb_gf4_mul_3_0_n59), .ZN(mult_lsb_gf4_mul_3_0_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_3_0_U8 ( .A(n113), .B(n117), .ZN(
        mult_lsb_gf4_mul_3_0_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_3_0_U7 ( .A(Y1_4xDP[0]), .B(Y1_4xDP[2]), .ZN(
        mult_lsb_gf4_mul_3_0_n61) );
  NAND2_X1 mult_lsb_gf4_mul_3_0_U6 ( .A1(mult_lsb_gf4_mul_3_0_n58), .A2(
        mult_lsb_gf4_mul_3_0_n60), .ZN(mult_lsb_gf4_mul_3_0_n55) );
  XOR2_X1 mult_lsb_gf4_mul_3_0_U5 ( .A(Y1_4xDP[1]), .B(Y1_4xDP[3]), .Z(
        mult_lsb_gf4_mul_3_0_n60) );
  XOR2_X1 mult_lsb_gf4_mul_3_0_U4 ( .A(n115), .B(n119), .Z(
        mult_lsb_gf4_mul_3_0_n58) );
  NOR2_X1 mult_lsb_gf4_mul_3_0_U3 ( .A1(mult_lsb_gf4_mul_3_0_n54), .A2(
        mult_lsb_gf4_mul_3_0_n53), .ZN(mult_lsb_gf4_mul_3_0_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_3_0_U2 ( .A(n113), .B(n115), .ZN(
        mult_lsb_gf4_mul_3_0_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_3_0_U1 ( .A(Y1_4xDP[0]), .B(Y1_4xDP[1]), .ZN(
        mult_lsb_gf4_mul_3_0_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_2_3_U29 ( .A(mult_lsb_gf4_mul_2_3_n77), .B(
        mult_lsb_gf4_mul_2_3_n76), .ZN(mult_lsb_Xi_mul_Yj_11__3_) );
  NAND2_X1 mult_lsb_gf4_mul_2_3_U28 ( .A1(n111), .A2(Y1_4xDP[15]), .ZN(
        mult_lsb_gf4_mul_2_3_n76) );
  XOR2_X1 mult_lsb_gf4_mul_2_3_U27 ( .A(mult_lsb_gf4_mul_2_3_n75), .B(
        mult_lsb_gf4_mul_2_3_n74), .Z(mult_lsb_gf4_mul_2_3_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_2_3_U26 ( .A(mult_lsb_gf4_mul_2_3_n73), .B(
        mult_lsb_gf4_mul_2_3_n72), .ZN(mult_lsb_Xi_mul_Yj_11__2_) );
  NAND2_X1 mult_lsb_gf4_mul_2_3_U25 ( .A1(n109), .A2(Y1_4xDP[14]), .ZN(
        mult_lsb_gf4_mul_2_3_n72) );
  XOR2_X1 mult_lsb_gf4_mul_2_3_U24 ( .A(mult_lsb_gf4_mul_2_3_n74), .B(
        mult_lsb_gf4_mul_2_3_n71), .Z(mult_lsb_gf4_mul_2_3_n73) );
  NOR2_X1 mult_lsb_gf4_mul_2_3_U23 ( .A1(mult_lsb_gf4_mul_2_3_n70), .A2(
        mult_lsb_gf4_mul_2_3_n69), .ZN(mult_lsb_gf4_mul_2_3_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_2_3_U22 ( .A(n109), .B(n111), .ZN(
        mult_lsb_gf4_mul_2_3_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_2_3_U21 ( .A(Y1_4xDP[14]), .B(Y1_4xDP[15]), .ZN(
        mult_lsb_gf4_mul_2_3_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_2_3_U20 ( .A(mult_lsb_gf4_mul_2_3_n68), .B(
        mult_lsb_gf4_mul_2_3_n67), .ZN(mult_lsb_Xi_mul_Yj_11__1_) );
  NAND2_X1 mult_lsb_gf4_mul_2_3_U19 ( .A1(n107), .A2(Y1_4xDP[13]), .ZN(
        mult_lsb_gf4_mul_2_3_n67) );
  XOR2_X1 mult_lsb_gf4_mul_2_3_U18 ( .A(mult_lsb_gf4_mul_2_3_n75), .B(
        mult_lsb_gf4_mul_2_3_n66), .Z(mult_lsb_gf4_mul_2_3_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_2_3_U17 ( .A(mult_lsb_gf4_mul_2_3_n65), .B(
        mult_lsb_gf4_mul_2_3_n64), .ZN(mult_lsb_gf4_mul_2_3_n75) );
  NAND2_X1 mult_lsb_gf4_mul_2_3_U16 ( .A1(mult_lsb_gf4_mul_2_3_n63), .A2(
        mult_lsb_gf4_mul_2_3_n62), .ZN(mult_lsb_gf4_mul_2_3_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_2_3_U15 ( .A(mult_lsb_gf4_mul_2_3_n61), .B(
        mult_lsb_gf4_mul_2_3_n60), .ZN(mult_lsb_gf4_mul_2_3_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_2_3_U14 ( .A(mult_lsb_gf4_mul_2_3_n59), .B(
        mult_lsb_gf4_mul_2_3_n58), .ZN(mult_lsb_gf4_mul_2_3_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_2_3_U13 ( .A(mult_lsb_gf4_mul_2_3_n57), .B(
        mult_lsb_gf4_mul_2_3_n56), .ZN(mult_lsb_Xi_mul_Yj_11__0_) );
  NAND2_X1 mult_lsb_gf4_mul_2_3_U12 ( .A1(n105), .A2(Y1_4xDP[12]), .ZN(
        mult_lsb_gf4_mul_2_3_n56) );
  XOR2_X1 mult_lsb_gf4_mul_2_3_U11 ( .A(mult_lsb_gf4_mul_2_3_n66), .B(
        mult_lsb_gf4_mul_2_3_n71), .Z(mult_lsb_gf4_mul_2_3_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_2_3_U10 ( .A(mult_lsb_gf4_mul_2_3_n55), .B(
        mult_lsb_gf4_mul_2_3_n65), .ZN(mult_lsb_gf4_mul_2_3_n71) );
  NOR2_X1 mult_lsb_gf4_mul_2_3_U9 ( .A1(mult_lsb_gf4_mul_2_3_n61), .A2(
        mult_lsb_gf4_mul_2_3_n59), .ZN(mult_lsb_gf4_mul_2_3_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_2_3_U8 ( .A(n105), .B(n109), .ZN(
        mult_lsb_gf4_mul_2_3_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_2_3_U7 ( .A(Y1_4xDP[12]), .B(Y1_4xDP[14]), .ZN(
        mult_lsb_gf4_mul_2_3_n61) );
  NAND2_X1 mult_lsb_gf4_mul_2_3_U6 ( .A1(mult_lsb_gf4_mul_2_3_n58), .A2(
        mult_lsb_gf4_mul_2_3_n60), .ZN(mult_lsb_gf4_mul_2_3_n55) );
  XOR2_X1 mult_lsb_gf4_mul_2_3_U5 ( .A(Y1_4xDP[13]), .B(Y1_4xDP[15]), .Z(
        mult_lsb_gf4_mul_2_3_n60) );
  XOR2_X1 mult_lsb_gf4_mul_2_3_U4 ( .A(n107), .B(n111), .Z(
        mult_lsb_gf4_mul_2_3_n58) );
  NOR2_X1 mult_lsb_gf4_mul_2_3_U3 ( .A1(mult_lsb_gf4_mul_2_3_n54), .A2(
        mult_lsb_gf4_mul_2_3_n53), .ZN(mult_lsb_gf4_mul_2_3_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_2_3_U2 ( .A(n105), .B(n107), .ZN(
        mult_lsb_gf4_mul_2_3_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_2_3_U1 ( .A(Y1_4xDP[12]), .B(Y1_4xDP[13]), .ZN(
        mult_lsb_gf4_mul_2_3_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U29 ( .A(mult_lsb_gf4_mul_2_2_n77), .B(
        mult_lsb_gf4_mul_2_2_n76), .ZN(mult_lsb_FFxDN[43]) );
  NAND2_X1 mult_lsb_gf4_mul_2_2_U28 ( .A1(n111), .A2(Y1_4xDP[11]), .ZN(
        mult_lsb_gf4_mul_2_2_n76) );
  XOR2_X1 mult_lsb_gf4_mul_2_2_U27 ( .A(mult_lsb_gf4_mul_2_2_n75), .B(
        mult_lsb_gf4_mul_2_2_n74), .Z(mult_lsb_gf4_mul_2_2_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U26 ( .A(mult_lsb_gf4_mul_2_2_n73), .B(
        mult_lsb_gf4_mul_2_2_n72), .ZN(mult_lsb_FFxDN[42]) );
  NAND2_X1 mult_lsb_gf4_mul_2_2_U25 ( .A1(n109), .A2(Y1_4xDP[10]), .ZN(
        mult_lsb_gf4_mul_2_2_n72) );
  XOR2_X1 mult_lsb_gf4_mul_2_2_U24 ( .A(mult_lsb_gf4_mul_2_2_n74), .B(
        mult_lsb_gf4_mul_2_2_n71), .Z(mult_lsb_gf4_mul_2_2_n73) );
  NOR2_X1 mult_lsb_gf4_mul_2_2_U23 ( .A1(mult_lsb_gf4_mul_2_2_n70), .A2(
        mult_lsb_gf4_mul_2_2_n69), .ZN(mult_lsb_gf4_mul_2_2_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U22 ( .A(n109), .B(n111), .ZN(
        mult_lsb_gf4_mul_2_2_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U21 ( .A(Y1_4xDP[10]), .B(Y1_4xDP[11]), .ZN(
        mult_lsb_gf4_mul_2_2_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U20 ( .A(mult_lsb_gf4_mul_2_2_n68), .B(
        mult_lsb_gf4_mul_2_2_n67), .ZN(mult_lsb_FFxDN[41]) );
  NAND2_X1 mult_lsb_gf4_mul_2_2_U19 ( .A1(n107), .A2(Y1_4xDP[9]), .ZN(
        mult_lsb_gf4_mul_2_2_n67) );
  XOR2_X1 mult_lsb_gf4_mul_2_2_U18 ( .A(mult_lsb_gf4_mul_2_2_n75), .B(
        mult_lsb_gf4_mul_2_2_n66), .Z(mult_lsb_gf4_mul_2_2_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U17 ( .A(mult_lsb_gf4_mul_2_2_n65), .B(
        mult_lsb_gf4_mul_2_2_n64), .ZN(mult_lsb_gf4_mul_2_2_n75) );
  NAND2_X1 mult_lsb_gf4_mul_2_2_U16 ( .A1(mult_lsb_gf4_mul_2_2_n63), .A2(
        mult_lsb_gf4_mul_2_2_n62), .ZN(mult_lsb_gf4_mul_2_2_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U15 ( .A(mult_lsb_gf4_mul_2_2_n61), .B(
        mult_lsb_gf4_mul_2_2_n60), .ZN(mult_lsb_gf4_mul_2_2_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U14 ( .A(mult_lsb_gf4_mul_2_2_n59), .B(
        mult_lsb_gf4_mul_2_2_n58), .ZN(mult_lsb_gf4_mul_2_2_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U13 ( .A(mult_lsb_gf4_mul_2_2_n57), .B(
        mult_lsb_gf4_mul_2_2_n56), .ZN(mult_lsb_FFxDN[40]) );
  NAND2_X1 mult_lsb_gf4_mul_2_2_U12 ( .A1(n105), .A2(Y1_4xDP[8]), .ZN(
        mult_lsb_gf4_mul_2_2_n56) );
  XOR2_X1 mult_lsb_gf4_mul_2_2_U11 ( .A(mult_lsb_gf4_mul_2_2_n66), .B(
        mult_lsb_gf4_mul_2_2_n71), .Z(mult_lsb_gf4_mul_2_2_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U10 ( .A(mult_lsb_gf4_mul_2_2_n55), .B(
        mult_lsb_gf4_mul_2_2_n65), .ZN(mult_lsb_gf4_mul_2_2_n71) );
  NOR2_X1 mult_lsb_gf4_mul_2_2_U9 ( .A1(mult_lsb_gf4_mul_2_2_n61), .A2(
        mult_lsb_gf4_mul_2_2_n59), .ZN(mult_lsb_gf4_mul_2_2_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U8 ( .A(n105), .B(n109), .ZN(
        mult_lsb_gf4_mul_2_2_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U7 ( .A(Y1_4xDP[8]), .B(Y1_4xDP[10]), .ZN(
        mult_lsb_gf4_mul_2_2_n61) );
  NAND2_X1 mult_lsb_gf4_mul_2_2_U6 ( .A1(mult_lsb_gf4_mul_2_2_n58), .A2(
        mult_lsb_gf4_mul_2_2_n60), .ZN(mult_lsb_gf4_mul_2_2_n55) );
  XOR2_X1 mult_lsb_gf4_mul_2_2_U5 ( .A(Y1_4xDP[9]), .B(Y1_4xDP[11]), .Z(
        mult_lsb_gf4_mul_2_2_n60) );
  XOR2_X1 mult_lsb_gf4_mul_2_2_U4 ( .A(n107), .B(n111), .Z(
        mult_lsb_gf4_mul_2_2_n58) );
  NOR2_X1 mult_lsb_gf4_mul_2_2_U3 ( .A1(mult_lsb_gf4_mul_2_2_n54), .A2(
        mult_lsb_gf4_mul_2_2_n53), .ZN(mult_lsb_gf4_mul_2_2_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U2 ( .A(n105), .B(n107), .ZN(
        mult_lsb_gf4_mul_2_2_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_2_2_U1 ( .A(Y1_4xDP[8]), .B(Y1_4xDP[9]), .ZN(
        mult_lsb_gf4_mul_2_2_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U29 ( .A(mult_lsb_gf4_mul_2_1_n77), .B(
        mult_lsb_gf4_mul_2_1_n76), .ZN(mult_lsb_Xi_mul_Yj_9__3_) );
  NAND2_X1 mult_lsb_gf4_mul_2_1_U28 ( .A1(n111), .A2(Y1_4xDP[7]), .ZN(
        mult_lsb_gf4_mul_2_1_n76) );
  XOR2_X1 mult_lsb_gf4_mul_2_1_U27 ( .A(mult_lsb_gf4_mul_2_1_n75), .B(
        mult_lsb_gf4_mul_2_1_n74), .Z(mult_lsb_gf4_mul_2_1_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U26 ( .A(mult_lsb_gf4_mul_2_1_n73), .B(
        mult_lsb_gf4_mul_2_1_n72), .ZN(mult_lsb_Xi_mul_Yj_9__2_) );
  NAND2_X1 mult_lsb_gf4_mul_2_1_U25 ( .A1(n109), .A2(Y1_4xDP[6]), .ZN(
        mult_lsb_gf4_mul_2_1_n72) );
  XOR2_X1 mult_lsb_gf4_mul_2_1_U24 ( .A(mult_lsb_gf4_mul_2_1_n74), .B(
        mult_lsb_gf4_mul_2_1_n71), .Z(mult_lsb_gf4_mul_2_1_n73) );
  NOR2_X1 mult_lsb_gf4_mul_2_1_U23 ( .A1(mult_lsb_gf4_mul_2_1_n70), .A2(
        mult_lsb_gf4_mul_2_1_n69), .ZN(mult_lsb_gf4_mul_2_1_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U22 ( .A(n109), .B(n111), .ZN(
        mult_lsb_gf4_mul_2_1_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U21 ( .A(Y1_4xDP[6]), .B(Y1_4xDP[7]), .ZN(
        mult_lsb_gf4_mul_2_1_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U20 ( .A(mult_lsb_gf4_mul_2_1_n68), .B(
        mult_lsb_gf4_mul_2_1_n67), .ZN(mult_lsb_Xi_mul_Yj_9__1_) );
  NAND2_X1 mult_lsb_gf4_mul_2_1_U19 ( .A1(n107), .A2(Y1_4xDP[5]), .ZN(
        mult_lsb_gf4_mul_2_1_n67) );
  XOR2_X1 mult_lsb_gf4_mul_2_1_U18 ( .A(mult_lsb_gf4_mul_2_1_n75), .B(
        mult_lsb_gf4_mul_2_1_n66), .Z(mult_lsb_gf4_mul_2_1_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U17 ( .A(mult_lsb_gf4_mul_2_1_n65), .B(
        mult_lsb_gf4_mul_2_1_n64), .ZN(mult_lsb_gf4_mul_2_1_n75) );
  NAND2_X1 mult_lsb_gf4_mul_2_1_U16 ( .A1(mult_lsb_gf4_mul_2_1_n63), .A2(
        mult_lsb_gf4_mul_2_1_n62), .ZN(mult_lsb_gf4_mul_2_1_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U15 ( .A(mult_lsb_gf4_mul_2_1_n61), .B(
        mult_lsb_gf4_mul_2_1_n60), .ZN(mult_lsb_gf4_mul_2_1_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U14 ( .A(mult_lsb_gf4_mul_2_1_n59), .B(
        mult_lsb_gf4_mul_2_1_n58), .ZN(mult_lsb_gf4_mul_2_1_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U13 ( .A(mult_lsb_gf4_mul_2_1_n57), .B(
        mult_lsb_gf4_mul_2_1_n56), .ZN(mult_lsb_Xi_mul_Yj_9__0_) );
  NAND2_X1 mult_lsb_gf4_mul_2_1_U12 ( .A1(n105), .A2(Y1_4xDP[4]), .ZN(
        mult_lsb_gf4_mul_2_1_n56) );
  XOR2_X1 mult_lsb_gf4_mul_2_1_U11 ( .A(mult_lsb_gf4_mul_2_1_n66), .B(
        mult_lsb_gf4_mul_2_1_n71), .Z(mult_lsb_gf4_mul_2_1_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U10 ( .A(mult_lsb_gf4_mul_2_1_n55), .B(
        mult_lsb_gf4_mul_2_1_n65), .ZN(mult_lsb_gf4_mul_2_1_n71) );
  NOR2_X1 mult_lsb_gf4_mul_2_1_U9 ( .A1(mult_lsb_gf4_mul_2_1_n61), .A2(
        mult_lsb_gf4_mul_2_1_n59), .ZN(mult_lsb_gf4_mul_2_1_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U8 ( .A(n105), .B(n109), .ZN(
        mult_lsb_gf4_mul_2_1_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U7 ( .A(Y1_4xDP[4]), .B(Y1_4xDP[6]), .ZN(
        mult_lsb_gf4_mul_2_1_n61) );
  NAND2_X1 mult_lsb_gf4_mul_2_1_U6 ( .A1(mult_lsb_gf4_mul_2_1_n58), .A2(
        mult_lsb_gf4_mul_2_1_n60), .ZN(mult_lsb_gf4_mul_2_1_n55) );
  XOR2_X1 mult_lsb_gf4_mul_2_1_U5 ( .A(Y1_4xDP[5]), .B(Y1_4xDP[7]), .Z(
        mult_lsb_gf4_mul_2_1_n60) );
  XOR2_X1 mult_lsb_gf4_mul_2_1_U4 ( .A(n107), .B(n111), .Z(
        mult_lsb_gf4_mul_2_1_n58) );
  NOR2_X1 mult_lsb_gf4_mul_2_1_U3 ( .A1(mult_lsb_gf4_mul_2_1_n54), .A2(
        mult_lsb_gf4_mul_2_1_n53), .ZN(mult_lsb_gf4_mul_2_1_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U2 ( .A(n105), .B(n107), .ZN(
        mult_lsb_gf4_mul_2_1_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_2_1_U1 ( .A(Y1_4xDP[4]), .B(Y1_4xDP[5]), .ZN(
        mult_lsb_gf4_mul_2_1_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U29 ( .A(mult_lsb_gf4_mul_2_0_n77), .B(
        mult_lsb_gf4_mul_2_0_n76), .ZN(mult_lsb_Xi_mul_Yj_8__3_) );
  NAND2_X1 mult_lsb_gf4_mul_2_0_U28 ( .A1(n111), .A2(Y1_4xDP[3]), .ZN(
        mult_lsb_gf4_mul_2_0_n76) );
  XOR2_X1 mult_lsb_gf4_mul_2_0_U27 ( .A(mult_lsb_gf4_mul_2_0_n75), .B(
        mult_lsb_gf4_mul_2_0_n74), .Z(mult_lsb_gf4_mul_2_0_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U26 ( .A(mult_lsb_gf4_mul_2_0_n73), .B(
        mult_lsb_gf4_mul_2_0_n72), .ZN(mult_lsb_Xi_mul_Yj_8__2_) );
  NAND2_X1 mult_lsb_gf4_mul_2_0_U25 ( .A1(n109), .A2(Y1_4xDP[2]), .ZN(
        mult_lsb_gf4_mul_2_0_n72) );
  XOR2_X1 mult_lsb_gf4_mul_2_0_U24 ( .A(mult_lsb_gf4_mul_2_0_n74), .B(
        mult_lsb_gf4_mul_2_0_n71), .Z(mult_lsb_gf4_mul_2_0_n73) );
  NOR2_X1 mult_lsb_gf4_mul_2_0_U23 ( .A1(mult_lsb_gf4_mul_2_0_n70), .A2(
        mult_lsb_gf4_mul_2_0_n69), .ZN(mult_lsb_gf4_mul_2_0_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U22 ( .A(n109), .B(n111), .ZN(
        mult_lsb_gf4_mul_2_0_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U21 ( .A(Y1_4xDP[2]), .B(Y1_4xDP[3]), .ZN(
        mult_lsb_gf4_mul_2_0_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U20 ( .A(mult_lsb_gf4_mul_2_0_n68), .B(
        mult_lsb_gf4_mul_2_0_n67), .ZN(mult_lsb_Xi_mul_Yj_8__1_) );
  NAND2_X1 mult_lsb_gf4_mul_2_0_U19 ( .A1(n107), .A2(Y1_4xDP[1]), .ZN(
        mult_lsb_gf4_mul_2_0_n67) );
  XOR2_X1 mult_lsb_gf4_mul_2_0_U18 ( .A(mult_lsb_gf4_mul_2_0_n75), .B(
        mult_lsb_gf4_mul_2_0_n66), .Z(mult_lsb_gf4_mul_2_0_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U17 ( .A(mult_lsb_gf4_mul_2_0_n65), .B(
        mult_lsb_gf4_mul_2_0_n64), .ZN(mult_lsb_gf4_mul_2_0_n75) );
  NAND2_X1 mult_lsb_gf4_mul_2_0_U16 ( .A1(mult_lsb_gf4_mul_2_0_n63), .A2(
        mult_lsb_gf4_mul_2_0_n62), .ZN(mult_lsb_gf4_mul_2_0_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U15 ( .A(mult_lsb_gf4_mul_2_0_n61), .B(
        mult_lsb_gf4_mul_2_0_n60), .ZN(mult_lsb_gf4_mul_2_0_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U14 ( .A(mult_lsb_gf4_mul_2_0_n59), .B(
        mult_lsb_gf4_mul_2_0_n58), .ZN(mult_lsb_gf4_mul_2_0_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U13 ( .A(mult_lsb_gf4_mul_2_0_n57), .B(
        mult_lsb_gf4_mul_2_0_n56), .ZN(mult_lsb_Xi_mul_Yj_8__0_) );
  NAND2_X1 mult_lsb_gf4_mul_2_0_U12 ( .A1(n105), .A2(Y1_4xDP[0]), .ZN(
        mult_lsb_gf4_mul_2_0_n56) );
  XOR2_X1 mult_lsb_gf4_mul_2_0_U11 ( .A(mult_lsb_gf4_mul_2_0_n66), .B(
        mult_lsb_gf4_mul_2_0_n71), .Z(mult_lsb_gf4_mul_2_0_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U10 ( .A(mult_lsb_gf4_mul_2_0_n55), .B(
        mult_lsb_gf4_mul_2_0_n65), .ZN(mult_lsb_gf4_mul_2_0_n71) );
  NOR2_X1 mult_lsb_gf4_mul_2_0_U9 ( .A1(mult_lsb_gf4_mul_2_0_n61), .A2(
        mult_lsb_gf4_mul_2_0_n59), .ZN(mult_lsb_gf4_mul_2_0_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U8 ( .A(n105), .B(n109), .ZN(
        mult_lsb_gf4_mul_2_0_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U7 ( .A(Y1_4xDP[0]), .B(Y1_4xDP[2]), .ZN(
        mult_lsb_gf4_mul_2_0_n61) );
  NAND2_X1 mult_lsb_gf4_mul_2_0_U6 ( .A1(mult_lsb_gf4_mul_2_0_n58), .A2(
        mult_lsb_gf4_mul_2_0_n60), .ZN(mult_lsb_gf4_mul_2_0_n55) );
  XOR2_X1 mult_lsb_gf4_mul_2_0_U5 ( .A(Y1_4xDP[1]), .B(Y1_4xDP[3]), .Z(
        mult_lsb_gf4_mul_2_0_n60) );
  XOR2_X1 mult_lsb_gf4_mul_2_0_U4 ( .A(n107), .B(n111), .Z(
        mult_lsb_gf4_mul_2_0_n58) );
  NOR2_X1 mult_lsb_gf4_mul_2_0_U3 ( .A1(mult_lsb_gf4_mul_2_0_n54), .A2(
        mult_lsb_gf4_mul_2_0_n53), .ZN(mult_lsb_gf4_mul_2_0_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U2 ( .A(n105), .B(n107), .ZN(
        mult_lsb_gf4_mul_2_0_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_2_0_U1 ( .A(Y1_4xDP[0]), .B(Y1_4xDP[1]), .ZN(
        mult_lsb_gf4_mul_2_0_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_1_3_U29 ( .A(mult_lsb_gf4_mul_1_3_n77), .B(
        mult_lsb_gf4_mul_1_3_n76), .ZN(mult_lsb_Xi_mul_Yj_7__3_) );
  NAND2_X1 mult_lsb_gf4_mul_1_3_U28 ( .A1(n103), .A2(Y1_4xDP[15]), .ZN(
        mult_lsb_gf4_mul_1_3_n76) );
  XOR2_X1 mult_lsb_gf4_mul_1_3_U27 ( .A(mult_lsb_gf4_mul_1_3_n75), .B(
        mult_lsb_gf4_mul_1_3_n74), .Z(mult_lsb_gf4_mul_1_3_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_1_3_U26 ( .A(mult_lsb_gf4_mul_1_3_n73), .B(
        mult_lsb_gf4_mul_1_3_n72), .ZN(mult_lsb_Xi_mul_Yj_7__2_) );
  NAND2_X1 mult_lsb_gf4_mul_1_3_U25 ( .A1(n101), .A2(Y1_4xDP[14]), .ZN(
        mult_lsb_gf4_mul_1_3_n72) );
  XOR2_X1 mult_lsb_gf4_mul_1_3_U24 ( .A(mult_lsb_gf4_mul_1_3_n74), .B(
        mult_lsb_gf4_mul_1_3_n71), .Z(mult_lsb_gf4_mul_1_3_n73) );
  NOR2_X1 mult_lsb_gf4_mul_1_3_U23 ( .A1(mult_lsb_gf4_mul_1_3_n70), .A2(
        mult_lsb_gf4_mul_1_3_n69), .ZN(mult_lsb_gf4_mul_1_3_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_1_3_U22 ( .A(n101), .B(n103), .ZN(
        mult_lsb_gf4_mul_1_3_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_1_3_U21 ( .A(Y1_4xDP[14]), .B(Y1_4xDP[15]), .ZN(
        mult_lsb_gf4_mul_1_3_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_1_3_U20 ( .A(mult_lsb_gf4_mul_1_3_n68), .B(
        mult_lsb_gf4_mul_1_3_n67), .ZN(mult_lsb_Xi_mul_Yj_7__1_) );
  NAND2_X1 mult_lsb_gf4_mul_1_3_U19 ( .A1(n99), .A2(Y1_4xDP[13]), .ZN(
        mult_lsb_gf4_mul_1_3_n67) );
  XOR2_X1 mult_lsb_gf4_mul_1_3_U18 ( .A(mult_lsb_gf4_mul_1_3_n75), .B(
        mult_lsb_gf4_mul_1_3_n66), .Z(mult_lsb_gf4_mul_1_3_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_1_3_U17 ( .A(mult_lsb_gf4_mul_1_3_n65), .B(
        mult_lsb_gf4_mul_1_3_n64), .ZN(mult_lsb_gf4_mul_1_3_n75) );
  NAND2_X1 mult_lsb_gf4_mul_1_3_U16 ( .A1(mult_lsb_gf4_mul_1_3_n63), .A2(
        mult_lsb_gf4_mul_1_3_n62), .ZN(mult_lsb_gf4_mul_1_3_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_1_3_U15 ( .A(mult_lsb_gf4_mul_1_3_n61), .B(
        mult_lsb_gf4_mul_1_3_n60), .ZN(mult_lsb_gf4_mul_1_3_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_1_3_U14 ( .A(mult_lsb_gf4_mul_1_3_n59), .B(
        mult_lsb_gf4_mul_1_3_n58), .ZN(mult_lsb_gf4_mul_1_3_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_1_3_U13 ( .A(mult_lsb_gf4_mul_1_3_n57), .B(
        mult_lsb_gf4_mul_1_3_n56), .ZN(mult_lsb_Xi_mul_Yj_7__0_) );
  NAND2_X1 mult_lsb_gf4_mul_1_3_U12 ( .A1(n97), .A2(Y1_4xDP[12]), .ZN(
        mult_lsb_gf4_mul_1_3_n56) );
  XOR2_X1 mult_lsb_gf4_mul_1_3_U11 ( .A(mult_lsb_gf4_mul_1_3_n66), .B(
        mult_lsb_gf4_mul_1_3_n71), .Z(mult_lsb_gf4_mul_1_3_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_1_3_U10 ( .A(mult_lsb_gf4_mul_1_3_n55), .B(
        mult_lsb_gf4_mul_1_3_n65), .ZN(mult_lsb_gf4_mul_1_3_n71) );
  NOR2_X1 mult_lsb_gf4_mul_1_3_U9 ( .A1(mult_lsb_gf4_mul_1_3_n61), .A2(
        mult_lsb_gf4_mul_1_3_n59), .ZN(mult_lsb_gf4_mul_1_3_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_1_3_U8 ( .A(n97), .B(n101), .ZN(
        mult_lsb_gf4_mul_1_3_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_1_3_U7 ( .A(Y1_4xDP[12]), .B(Y1_4xDP[14]), .ZN(
        mult_lsb_gf4_mul_1_3_n61) );
  NAND2_X1 mult_lsb_gf4_mul_1_3_U6 ( .A1(mult_lsb_gf4_mul_1_3_n58), .A2(
        mult_lsb_gf4_mul_1_3_n60), .ZN(mult_lsb_gf4_mul_1_3_n55) );
  XOR2_X1 mult_lsb_gf4_mul_1_3_U5 ( .A(Y1_4xDP[13]), .B(Y1_4xDP[15]), .Z(
        mult_lsb_gf4_mul_1_3_n60) );
  XOR2_X1 mult_lsb_gf4_mul_1_3_U4 ( .A(n99), .B(n103), .Z(
        mult_lsb_gf4_mul_1_3_n58) );
  NOR2_X1 mult_lsb_gf4_mul_1_3_U3 ( .A1(mult_lsb_gf4_mul_1_3_n54), .A2(
        mult_lsb_gf4_mul_1_3_n53), .ZN(mult_lsb_gf4_mul_1_3_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_1_3_U2 ( .A(n97), .B(n99), .ZN(
        mult_lsb_gf4_mul_1_3_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_1_3_U1 ( .A(Y1_4xDP[12]), .B(Y1_4xDP[13]), .ZN(
        mult_lsb_gf4_mul_1_3_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U29 ( .A(mult_lsb_gf4_mul_1_2_n77), .B(
        mult_lsb_gf4_mul_1_2_n76), .ZN(mult_lsb_Xi_mul_Yj_6__3_) );
  NAND2_X1 mult_lsb_gf4_mul_1_2_U28 ( .A1(n103), .A2(Y1_4xDP[11]), .ZN(
        mult_lsb_gf4_mul_1_2_n76) );
  XOR2_X1 mult_lsb_gf4_mul_1_2_U27 ( .A(mult_lsb_gf4_mul_1_2_n75), .B(
        mult_lsb_gf4_mul_1_2_n74), .Z(mult_lsb_gf4_mul_1_2_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U26 ( .A(mult_lsb_gf4_mul_1_2_n73), .B(
        mult_lsb_gf4_mul_1_2_n72), .ZN(mult_lsb_Xi_mul_Yj_6__2_) );
  NAND2_X1 mult_lsb_gf4_mul_1_2_U25 ( .A1(n101), .A2(Y1_4xDP[10]), .ZN(
        mult_lsb_gf4_mul_1_2_n72) );
  XOR2_X1 mult_lsb_gf4_mul_1_2_U24 ( .A(mult_lsb_gf4_mul_1_2_n74), .B(
        mult_lsb_gf4_mul_1_2_n71), .Z(mult_lsb_gf4_mul_1_2_n73) );
  NOR2_X1 mult_lsb_gf4_mul_1_2_U23 ( .A1(mult_lsb_gf4_mul_1_2_n70), .A2(
        mult_lsb_gf4_mul_1_2_n69), .ZN(mult_lsb_gf4_mul_1_2_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U22 ( .A(n101), .B(n103), .ZN(
        mult_lsb_gf4_mul_1_2_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U21 ( .A(Y1_4xDP[10]), .B(Y1_4xDP[11]), .ZN(
        mult_lsb_gf4_mul_1_2_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U20 ( .A(mult_lsb_gf4_mul_1_2_n68), .B(
        mult_lsb_gf4_mul_1_2_n67), .ZN(mult_lsb_Xi_mul_Yj_6__1_) );
  NAND2_X1 mult_lsb_gf4_mul_1_2_U19 ( .A1(n99), .A2(Y1_4xDP[9]), .ZN(
        mult_lsb_gf4_mul_1_2_n67) );
  XOR2_X1 mult_lsb_gf4_mul_1_2_U18 ( .A(mult_lsb_gf4_mul_1_2_n75), .B(
        mult_lsb_gf4_mul_1_2_n66), .Z(mult_lsb_gf4_mul_1_2_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U17 ( .A(mult_lsb_gf4_mul_1_2_n65), .B(
        mult_lsb_gf4_mul_1_2_n64), .ZN(mult_lsb_gf4_mul_1_2_n75) );
  NAND2_X1 mult_lsb_gf4_mul_1_2_U16 ( .A1(mult_lsb_gf4_mul_1_2_n63), .A2(
        mult_lsb_gf4_mul_1_2_n62), .ZN(mult_lsb_gf4_mul_1_2_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U15 ( .A(mult_lsb_gf4_mul_1_2_n61), .B(
        mult_lsb_gf4_mul_1_2_n60), .ZN(mult_lsb_gf4_mul_1_2_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U14 ( .A(mult_lsb_gf4_mul_1_2_n59), .B(
        mult_lsb_gf4_mul_1_2_n58), .ZN(mult_lsb_gf4_mul_1_2_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U13 ( .A(mult_lsb_gf4_mul_1_2_n57), .B(
        mult_lsb_gf4_mul_1_2_n56), .ZN(mult_lsb_Xi_mul_Yj_6__0_) );
  NAND2_X1 mult_lsb_gf4_mul_1_2_U12 ( .A1(n97), .A2(Y1_4xDP[8]), .ZN(
        mult_lsb_gf4_mul_1_2_n56) );
  XOR2_X1 mult_lsb_gf4_mul_1_2_U11 ( .A(mult_lsb_gf4_mul_1_2_n66), .B(
        mult_lsb_gf4_mul_1_2_n71), .Z(mult_lsb_gf4_mul_1_2_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U10 ( .A(mult_lsb_gf4_mul_1_2_n55), .B(
        mult_lsb_gf4_mul_1_2_n65), .ZN(mult_lsb_gf4_mul_1_2_n71) );
  NOR2_X1 mult_lsb_gf4_mul_1_2_U9 ( .A1(mult_lsb_gf4_mul_1_2_n61), .A2(
        mult_lsb_gf4_mul_1_2_n59), .ZN(mult_lsb_gf4_mul_1_2_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U8 ( .A(n97), .B(n101), .ZN(
        mult_lsb_gf4_mul_1_2_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U7 ( .A(Y1_4xDP[8]), .B(Y1_4xDP[10]), .ZN(
        mult_lsb_gf4_mul_1_2_n61) );
  NAND2_X1 mult_lsb_gf4_mul_1_2_U6 ( .A1(mult_lsb_gf4_mul_1_2_n58), .A2(
        mult_lsb_gf4_mul_1_2_n60), .ZN(mult_lsb_gf4_mul_1_2_n55) );
  XOR2_X1 mult_lsb_gf4_mul_1_2_U5 ( .A(Y1_4xDP[9]), .B(Y1_4xDP[11]), .Z(
        mult_lsb_gf4_mul_1_2_n60) );
  XOR2_X1 mult_lsb_gf4_mul_1_2_U4 ( .A(n99), .B(n103), .Z(
        mult_lsb_gf4_mul_1_2_n58) );
  NOR2_X1 mult_lsb_gf4_mul_1_2_U3 ( .A1(mult_lsb_gf4_mul_1_2_n54), .A2(
        mult_lsb_gf4_mul_1_2_n53), .ZN(mult_lsb_gf4_mul_1_2_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U2 ( .A(n97), .B(n99), .ZN(
        mult_lsb_gf4_mul_1_2_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_1_2_U1 ( .A(Y1_4xDP[8]), .B(Y1_4xDP[9]), .ZN(
        mult_lsb_gf4_mul_1_2_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U29 ( .A(mult_lsb_gf4_mul_1_1_n77), .B(
        mult_lsb_gf4_mul_1_1_n76), .ZN(mult_lsb_FFxDN[23]) );
  NAND2_X1 mult_lsb_gf4_mul_1_1_U28 ( .A1(n103), .A2(Y1_4xDP[7]), .ZN(
        mult_lsb_gf4_mul_1_1_n76) );
  XOR2_X1 mult_lsb_gf4_mul_1_1_U27 ( .A(mult_lsb_gf4_mul_1_1_n75), .B(
        mult_lsb_gf4_mul_1_1_n74), .Z(mult_lsb_gf4_mul_1_1_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U26 ( .A(mult_lsb_gf4_mul_1_1_n73), .B(
        mult_lsb_gf4_mul_1_1_n72), .ZN(mult_lsb_FFxDN[22]) );
  NAND2_X1 mult_lsb_gf4_mul_1_1_U25 ( .A1(n101), .A2(Y1_4xDP[6]), .ZN(
        mult_lsb_gf4_mul_1_1_n72) );
  XOR2_X1 mult_lsb_gf4_mul_1_1_U24 ( .A(mult_lsb_gf4_mul_1_1_n74), .B(
        mult_lsb_gf4_mul_1_1_n71), .Z(mult_lsb_gf4_mul_1_1_n73) );
  NOR2_X1 mult_lsb_gf4_mul_1_1_U23 ( .A1(mult_lsb_gf4_mul_1_1_n70), .A2(
        mult_lsb_gf4_mul_1_1_n69), .ZN(mult_lsb_gf4_mul_1_1_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U22 ( .A(n101), .B(n103), .ZN(
        mult_lsb_gf4_mul_1_1_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U21 ( .A(Y1_4xDP[6]), .B(Y1_4xDP[7]), .ZN(
        mult_lsb_gf4_mul_1_1_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U20 ( .A(mult_lsb_gf4_mul_1_1_n68), .B(
        mult_lsb_gf4_mul_1_1_n67), .ZN(mult_lsb_FFxDN[21]) );
  NAND2_X1 mult_lsb_gf4_mul_1_1_U19 ( .A1(n99), .A2(Y1_4xDP[5]), .ZN(
        mult_lsb_gf4_mul_1_1_n67) );
  XOR2_X1 mult_lsb_gf4_mul_1_1_U18 ( .A(mult_lsb_gf4_mul_1_1_n75), .B(
        mult_lsb_gf4_mul_1_1_n66), .Z(mult_lsb_gf4_mul_1_1_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U17 ( .A(mult_lsb_gf4_mul_1_1_n65), .B(
        mult_lsb_gf4_mul_1_1_n64), .ZN(mult_lsb_gf4_mul_1_1_n75) );
  NAND2_X1 mult_lsb_gf4_mul_1_1_U16 ( .A1(mult_lsb_gf4_mul_1_1_n63), .A2(
        mult_lsb_gf4_mul_1_1_n62), .ZN(mult_lsb_gf4_mul_1_1_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U15 ( .A(mult_lsb_gf4_mul_1_1_n61), .B(
        mult_lsb_gf4_mul_1_1_n60), .ZN(mult_lsb_gf4_mul_1_1_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U14 ( .A(mult_lsb_gf4_mul_1_1_n59), .B(
        mult_lsb_gf4_mul_1_1_n58), .ZN(mult_lsb_gf4_mul_1_1_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U13 ( .A(mult_lsb_gf4_mul_1_1_n57), .B(
        mult_lsb_gf4_mul_1_1_n56), .ZN(mult_lsb_FFxDN[20]) );
  NAND2_X1 mult_lsb_gf4_mul_1_1_U12 ( .A1(n97), .A2(Y1_4xDP[4]), .ZN(
        mult_lsb_gf4_mul_1_1_n56) );
  XOR2_X1 mult_lsb_gf4_mul_1_1_U11 ( .A(mult_lsb_gf4_mul_1_1_n66), .B(
        mult_lsb_gf4_mul_1_1_n71), .Z(mult_lsb_gf4_mul_1_1_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U10 ( .A(mult_lsb_gf4_mul_1_1_n55), .B(
        mult_lsb_gf4_mul_1_1_n65), .ZN(mult_lsb_gf4_mul_1_1_n71) );
  NOR2_X1 mult_lsb_gf4_mul_1_1_U9 ( .A1(mult_lsb_gf4_mul_1_1_n61), .A2(
        mult_lsb_gf4_mul_1_1_n59), .ZN(mult_lsb_gf4_mul_1_1_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U8 ( .A(n97), .B(n101), .ZN(
        mult_lsb_gf4_mul_1_1_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U7 ( .A(Y1_4xDP[4]), .B(Y1_4xDP[6]), .ZN(
        mult_lsb_gf4_mul_1_1_n61) );
  NAND2_X1 mult_lsb_gf4_mul_1_1_U6 ( .A1(mult_lsb_gf4_mul_1_1_n58), .A2(
        mult_lsb_gf4_mul_1_1_n60), .ZN(mult_lsb_gf4_mul_1_1_n55) );
  XOR2_X1 mult_lsb_gf4_mul_1_1_U5 ( .A(Y1_4xDP[5]), .B(Y1_4xDP[7]), .Z(
        mult_lsb_gf4_mul_1_1_n60) );
  XOR2_X1 mult_lsb_gf4_mul_1_1_U4 ( .A(n99), .B(n103), .Z(
        mult_lsb_gf4_mul_1_1_n58) );
  NOR2_X1 mult_lsb_gf4_mul_1_1_U3 ( .A1(mult_lsb_gf4_mul_1_1_n54), .A2(
        mult_lsb_gf4_mul_1_1_n53), .ZN(mult_lsb_gf4_mul_1_1_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U2 ( .A(n97), .B(n99), .ZN(
        mult_lsb_gf4_mul_1_1_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_1_1_U1 ( .A(Y1_4xDP[4]), .B(Y1_4xDP[5]), .ZN(
        mult_lsb_gf4_mul_1_1_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U29 ( .A(mult_lsb_gf4_mul_1_0_n77), .B(
        mult_lsb_gf4_mul_1_0_n76), .ZN(mult_lsb_Xi_mul_Yj_4__3_) );
  NAND2_X1 mult_lsb_gf4_mul_1_0_U28 ( .A1(n103), .A2(Y1_4xDP[3]), .ZN(
        mult_lsb_gf4_mul_1_0_n76) );
  XOR2_X1 mult_lsb_gf4_mul_1_0_U27 ( .A(mult_lsb_gf4_mul_1_0_n75), .B(
        mult_lsb_gf4_mul_1_0_n74), .Z(mult_lsb_gf4_mul_1_0_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U26 ( .A(mult_lsb_gf4_mul_1_0_n73), .B(
        mult_lsb_gf4_mul_1_0_n72), .ZN(mult_lsb_Xi_mul_Yj_4__2_) );
  NAND2_X1 mult_lsb_gf4_mul_1_0_U25 ( .A1(n101), .A2(Y1_4xDP[2]), .ZN(
        mult_lsb_gf4_mul_1_0_n72) );
  XOR2_X1 mult_lsb_gf4_mul_1_0_U24 ( .A(mult_lsb_gf4_mul_1_0_n74), .B(
        mult_lsb_gf4_mul_1_0_n71), .Z(mult_lsb_gf4_mul_1_0_n73) );
  NOR2_X1 mult_lsb_gf4_mul_1_0_U23 ( .A1(mult_lsb_gf4_mul_1_0_n70), .A2(
        mult_lsb_gf4_mul_1_0_n69), .ZN(mult_lsb_gf4_mul_1_0_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U22 ( .A(n101), .B(n103), .ZN(
        mult_lsb_gf4_mul_1_0_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U21 ( .A(Y1_4xDP[2]), .B(Y1_4xDP[3]), .ZN(
        mult_lsb_gf4_mul_1_0_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U20 ( .A(mult_lsb_gf4_mul_1_0_n68), .B(
        mult_lsb_gf4_mul_1_0_n67), .ZN(mult_lsb_Xi_mul_Yj_4__1_) );
  NAND2_X1 mult_lsb_gf4_mul_1_0_U19 ( .A1(n99), .A2(Y1_4xDP[1]), .ZN(
        mult_lsb_gf4_mul_1_0_n67) );
  XOR2_X1 mult_lsb_gf4_mul_1_0_U18 ( .A(mult_lsb_gf4_mul_1_0_n75), .B(
        mult_lsb_gf4_mul_1_0_n66), .Z(mult_lsb_gf4_mul_1_0_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U17 ( .A(mult_lsb_gf4_mul_1_0_n65), .B(
        mult_lsb_gf4_mul_1_0_n64), .ZN(mult_lsb_gf4_mul_1_0_n75) );
  NAND2_X1 mult_lsb_gf4_mul_1_0_U16 ( .A1(mult_lsb_gf4_mul_1_0_n63), .A2(
        mult_lsb_gf4_mul_1_0_n62), .ZN(mult_lsb_gf4_mul_1_0_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U15 ( .A(mult_lsb_gf4_mul_1_0_n61), .B(
        mult_lsb_gf4_mul_1_0_n60), .ZN(mult_lsb_gf4_mul_1_0_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U14 ( .A(mult_lsb_gf4_mul_1_0_n59), .B(
        mult_lsb_gf4_mul_1_0_n58), .ZN(mult_lsb_gf4_mul_1_0_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U13 ( .A(mult_lsb_gf4_mul_1_0_n57), .B(
        mult_lsb_gf4_mul_1_0_n56), .ZN(mult_lsb_Xi_mul_Yj_4__0_) );
  NAND2_X1 mult_lsb_gf4_mul_1_0_U12 ( .A1(n97), .A2(Y1_4xDP[0]), .ZN(
        mult_lsb_gf4_mul_1_0_n56) );
  XOR2_X1 mult_lsb_gf4_mul_1_0_U11 ( .A(mult_lsb_gf4_mul_1_0_n66), .B(
        mult_lsb_gf4_mul_1_0_n71), .Z(mult_lsb_gf4_mul_1_0_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U10 ( .A(mult_lsb_gf4_mul_1_0_n55), .B(
        mult_lsb_gf4_mul_1_0_n65), .ZN(mult_lsb_gf4_mul_1_0_n71) );
  NOR2_X1 mult_lsb_gf4_mul_1_0_U9 ( .A1(mult_lsb_gf4_mul_1_0_n61), .A2(
        mult_lsb_gf4_mul_1_0_n59), .ZN(mult_lsb_gf4_mul_1_0_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U8 ( .A(n97), .B(n101), .ZN(
        mult_lsb_gf4_mul_1_0_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U7 ( .A(Y1_4xDP[0]), .B(Y1_4xDP[2]), .ZN(
        mult_lsb_gf4_mul_1_0_n61) );
  NAND2_X1 mult_lsb_gf4_mul_1_0_U6 ( .A1(mult_lsb_gf4_mul_1_0_n58), .A2(
        mult_lsb_gf4_mul_1_0_n60), .ZN(mult_lsb_gf4_mul_1_0_n55) );
  XOR2_X1 mult_lsb_gf4_mul_1_0_U5 ( .A(Y1_4xDP[1]), .B(Y1_4xDP[3]), .Z(
        mult_lsb_gf4_mul_1_0_n60) );
  XOR2_X1 mult_lsb_gf4_mul_1_0_U4 ( .A(n99), .B(n103), .Z(
        mult_lsb_gf4_mul_1_0_n58) );
  NOR2_X1 mult_lsb_gf4_mul_1_0_U3 ( .A1(mult_lsb_gf4_mul_1_0_n54), .A2(
        mult_lsb_gf4_mul_1_0_n53), .ZN(mult_lsb_gf4_mul_1_0_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U2 ( .A(n97), .B(n99), .ZN(
        mult_lsb_gf4_mul_1_0_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_1_0_U1 ( .A(Y1_4xDP[0]), .B(Y1_4xDP[1]), .ZN(
        mult_lsb_gf4_mul_1_0_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_0_3_U29 ( .A(mult_lsb_gf4_mul_0_3_n77), .B(
        mult_lsb_gf4_mul_0_3_n76), .ZN(mult_lsb_Xi_mul_Yj_3__3_) );
  NAND2_X1 mult_lsb_gf4_mul_0_3_U28 ( .A1(n95), .A2(Y1_4xDP[15]), .ZN(
        mult_lsb_gf4_mul_0_3_n76) );
  XOR2_X1 mult_lsb_gf4_mul_0_3_U27 ( .A(mult_lsb_gf4_mul_0_3_n75), .B(
        mult_lsb_gf4_mul_0_3_n74), .Z(mult_lsb_gf4_mul_0_3_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_0_3_U26 ( .A(mult_lsb_gf4_mul_0_3_n73), .B(
        mult_lsb_gf4_mul_0_3_n72), .ZN(mult_lsb_Xi_mul_Yj_3__2_) );
  NAND2_X1 mult_lsb_gf4_mul_0_3_U25 ( .A1(n93), .A2(Y1_4xDP[14]), .ZN(
        mult_lsb_gf4_mul_0_3_n72) );
  XOR2_X1 mult_lsb_gf4_mul_0_3_U24 ( .A(mult_lsb_gf4_mul_0_3_n74), .B(
        mult_lsb_gf4_mul_0_3_n71), .Z(mult_lsb_gf4_mul_0_3_n73) );
  NOR2_X1 mult_lsb_gf4_mul_0_3_U23 ( .A1(mult_lsb_gf4_mul_0_3_n70), .A2(
        mult_lsb_gf4_mul_0_3_n69), .ZN(mult_lsb_gf4_mul_0_3_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_0_3_U22 ( .A(n93), .B(n95), .ZN(
        mult_lsb_gf4_mul_0_3_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_0_3_U21 ( .A(Y1_4xDP[14]), .B(Y1_4xDP[15]), .ZN(
        mult_lsb_gf4_mul_0_3_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_0_3_U20 ( .A(mult_lsb_gf4_mul_0_3_n68), .B(
        mult_lsb_gf4_mul_0_3_n67), .ZN(mult_lsb_Xi_mul_Yj_3__1_) );
  NAND2_X1 mult_lsb_gf4_mul_0_3_U19 ( .A1(n91), .A2(Y1_4xDP[13]), .ZN(
        mult_lsb_gf4_mul_0_3_n67) );
  XOR2_X1 mult_lsb_gf4_mul_0_3_U18 ( .A(mult_lsb_gf4_mul_0_3_n75), .B(
        mult_lsb_gf4_mul_0_3_n66), .Z(mult_lsb_gf4_mul_0_3_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_0_3_U17 ( .A(mult_lsb_gf4_mul_0_3_n65), .B(
        mult_lsb_gf4_mul_0_3_n64), .ZN(mult_lsb_gf4_mul_0_3_n75) );
  NAND2_X1 mult_lsb_gf4_mul_0_3_U16 ( .A1(mult_lsb_gf4_mul_0_3_n63), .A2(
        mult_lsb_gf4_mul_0_3_n62), .ZN(mult_lsb_gf4_mul_0_3_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_0_3_U15 ( .A(mult_lsb_gf4_mul_0_3_n61), .B(
        mult_lsb_gf4_mul_0_3_n60), .ZN(mult_lsb_gf4_mul_0_3_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_0_3_U14 ( .A(mult_lsb_gf4_mul_0_3_n59), .B(
        mult_lsb_gf4_mul_0_3_n58), .ZN(mult_lsb_gf4_mul_0_3_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_0_3_U13 ( .A(mult_lsb_gf4_mul_0_3_n57), .B(
        mult_lsb_gf4_mul_0_3_n56), .ZN(mult_lsb_Xi_mul_Yj_3__0_) );
  NAND2_X1 mult_lsb_gf4_mul_0_3_U12 ( .A1(n89), .A2(Y1_4xDP[12]), .ZN(
        mult_lsb_gf4_mul_0_3_n56) );
  XOR2_X1 mult_lsb_gf4_mul_0_3_U11 ( .A(mult_lsb_gf4_mul_0_3_n66), .B(
        mult_lsb_gf4_mul_0_3_n71), .Z(mult_lsb_gf4_mul_0_3_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_0_3_U10 ( .A(mult_lsb_gf4_mul_0_3_n55), .B(
        mult_lsb_gf4_mul_0_3_n65), .ZN(mult_lsb_gf4_mul_0_3_n71) );
  NOR2_X1 mult_lsb_gf4_mul_0_3_U9 ( .A1(mult_lsb_gf4_mul_0_3_n61), .A2(
        mult_lsb_gf4_mul_0_3_n59), .ZN(mult_lsb_gf4_mul_0_3_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_0_3_U8 ( .A(n89), .B(n93), .ZN(
        mult_lsb_gf4_mul_0_3_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_0_3_U7 ( .A(Y1_4xDP[12]), .B(Y1_4xDP[14]), .ZN(
        mult_lsb_gf4_mul_0_3_n61) );
  NAND2_X1 mult_lsb_gf4_mul_0_3_U6 ( .A1(mult_lsb_gf4_mul_0_3_n58), .A2(
        mult_lsb_gf4_mul_0_3_n60), .ZN(mult_lsb_gf4_mul_0_3_n55) );
  XOR2_X1 mult_lsb_gf4_mul_0_3_U5 ( .A(Y1_4xDP[13]), .B(Y1_4xDP[15]), .Z(
        mult_lsb_gf4_mul_0_3_n60) );
  XOR2_X1 mult_lsb_gf4_mul_0_3_U4 ( .A(n91), .B(n95), .Z(
        mult_lsb_gf4_mul_0_3_n58) );
  NOR2_X1 mult_lsb_gf4_mul_0_3_U3 ( .A1(mult_lsb_gf4_mul_0_3_n54), .A2(
        mult_lsb_gf4_mul_0_3_n53), .ZN(mult_lsb_gf4_mul_0_3_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_0_3_U2 ( .A(n89), .B(n91), .ZN(
        mult_lsb_gf4_mul_0_3_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_0_3_U1 ( .A(Y1_4xDP[12]), .B(Y1_4xDP[13]), .ZN(
        mult_lsb_gf4_mul_0_3_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U29 ( .A(mult_lsb_gf4_mul_0_2_n77), .B(
        mult_lsb_gf4_mul_0_2_n76), .ZN(mult_lsb_Xi_mul_Yj_2__3_) );
  NAND2_X1 mult_lsb_gf4_mul_0_2_U28 ( .A1(n95), .A2(Y1_4xDP[11]), .ZN(
        mult_lsb_gf4_mul_0_2_n76) );
  XOR2_X1 mult_lsb_gf4_mul_0_2_U27 ( .A(mult_lsb_gf4_mul_0_2_n75), .B(
        mult_lsb_gf4_mul_0_2_n74), .Z(mult_lsb_gf4_mul_0_2_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U26 ( .A(mult_lsb_gf4_mul_0_2_n73), .B(
        mult_lsb_gf4_mul_0_2_n72), .ZN(mult_lsb_Xi_mul_Yj_2__2_) );
  NAND2_X1 mult_lsb_gf4_mul_0_2_U25 ( .A1(n93), .A2(Y1_4xDP[10]), .ZN(
        mult_lsb_gf4_mul_0_2_n72) );
  XOR2_X1 mult_lsb_gf4_mul_0_2_U24 ( .A(mult_lsb_gf4_mul_0_2_n74), .B(
        mult_lsb_gf4_mul_0_2_n71), .Z(mult_lsb_gf4_mul_0_2_n73) );
  NOR2_X1 mult_lsb_gf4_mul_0_2_U23 ( .A1(mult_lsb_gf4_mul_0_2_n70), .A2(
        mult_lsb_gf4_mul_0_2_n69), .ZN(mult_lsb_gf4_mul_0_2_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U22 ( .A(n93), .B(n95), .ZN(
        mult_lsb_gf4_mul_0_2_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U21 ( .A(Y1_4xDP[10]), .B(Y1_4xDP[11]), .ZN(
        mult_lsb_gf4_mul_0_2_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U20 ( .A(mult_lsb_gf4_mul_0_2_n68), .B(
        mult_lsb_gf4_mul_0_2_n67), .ZN(mult_lsb_Xi_mul_Yj_2__1_) );
  NAND2_X1 mult_lsb_gf4_mul_0_2_U19 ( .A1(n91), .A2(Y1_4xDP[9]), .ZN(
        mult_lsb_gf4_mul_0_2_n67) );
  XOR2_X1 mult_lsb_gf4_mul_0_2_U18 ( .A(mult_lsb_gf4_mul_0_2_n75), .B(
        mult_lsb_gf4_mul_0_2_n66), .Z(mult_lsb_gf4_mul_0_2_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U17 ( .A(mult_lsb_gf4_mul_0_2_n65), .B(
        mult_lsb_gf4_mul_0_2_n64), .ZN(mult_lsb_gf4_mul_0_2_n75) );
  NAND2_X1 mult_lsb_gf4_mul_0_2_U16 ( .A1(mult_lsb_gf4_mul_0_2_n63), .A2(
        mult_lsb_gf4_mul_0_2_n62), .ZN(mult_lsb_gf4_mul_0_2_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U15 ( .A(mult_lsb_gf4_mul_0_2_n61), .B(
        mult_lsb_gf4_mul_0_2_n60), .ZN(mult_lsb_gf4_mul_0_2_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U14 ( .A(mult_lsb_gf4_mul_0_2_n59), .B(
        mult_lsb_gf4_mul_0_2_n58), .ZN(mult_lsb_gf4_mul_0_2_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U13 ( .A(mult_lsb_gf4_mul_0_2_n57), .B(
        mult_lsb_gf4_mul_0_2_n56), .ZN(mult_lsb_Xi_mul_Yj_2__0_) );
  NAND2_X1 mult_lsb_gf4_mul_0_2_U12 ( .A1(n89), .A2(Y1_4xDP[8]), .ZN(
        mult_lsb_gf4_mul_0_2_n56) );
  XOR2_X1 mult_lsb_gf4_mul_0_2_U11 ( .A(mult_lsb_gf4_mul_0_2_n66), .B(
        mult_lsb_gf4_mul_0_2_n71), .Z(mult_lsb_gf4_mul_0_2_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U10 ( .A(mult_lsb_gf4_mul_0_2_n55), .B(
        mult_lsb_gf4_mul_0_2_n65), .ZN(mult_lsb_gf4_mul_0_2_n71) );
  NOR2_X1 mult_lsb_gf4_mul_0_2_U9 ( .A1(mult_lsb_gf4_mul_0_2_n61), .A2(
        mult_lsb_gf4_mul_0_2_n59), .ZN(mult_lsb_gf4_mul_0_2_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U8 ( .A(n89), .B(n93), .ZN(
        mult_lsb_gf4_mul_0_2_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U7 ( .A(Y1_4xDP[8]), .B(Y1_4xDP[10]), .ZN(
        mult_lsb_gf4_mul_0_2_n61) );
  NAND2_X1 mult_lsb_gf4_mul_0_2_U6 ( .A1(mult_lsb_gf4_mul_0_2_n58), .A2(
        mult_lsb_gf4_mul_0_2_n60), .ZN(mult_lsb_gf4_mul_0_2_n55) );
  XOR2_X1 mult_lsb_gf4_mul_0_2_U5 ( .A(Y1_4xDP[9]), .B(Y1_4xDP[11]), .Z(
        mult_lsb_gf4_mul_0_2_n60) );
  XOR2_X1 mult_lsb_gf4_mul_0_2_U4 ( .A(n91), .B(n95), .Z(
        mult_lsb_gf4_mul_0_2_n58) );
  NOR2_X1 mult_lsb_gf4_mul_0_2_U3 ( .A1(mult_lsb_gf4_mul_0_2_n54), .A2(
        mult_lsb_gf4_mul_0_2_n53), .ZN(mult_lsb_gf4_mul_0_2_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U2 ( .A(n89), .B(n91), .ZN(
        mult_lsb_gf4_mul_0_2_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_0_2_U1 ( .A(Y1_4xDP[8]), .B(Y1_4xDP[9]), .ZN(
        mult_lsb_gf4_mul_0_2_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U29 ( .A(mult_lsb_gf4_mul_0_1_n77), .B(
        mult_lsb_gf4_mul_0_1_n76), .ZN(mult_lsb_Xi_mul_Yj_1__3_) );
  NAND2_X1 mult_lsb_gf4_mul_0_1_U28 ( .A1(n95), .A2(Y1_4xDP[7]), .ZN(
        mult_lsb_gf4_mul_0_1_n76) );
  XOR2_X1 mult_lsb_gf4_mul_0_1_U27 ( .A(mult_lsb_gf4_mul_0_1_n75), .B(
        mult_lsb_gf4_mul_0_1_n74), .Z(mult_lsb_gf4_mul_0_1_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U26 ( .A(mult_lsb_gf4_mul_0_1_n73), .B(
        mult_lsb_gf4_mul_0_1_n72), .ZN(mult_lsb_Xi_mul_Yj_1__2_) );
  NAND2_X1 mult_lsb_gf4_mul_0_1_U25 ( .A1(n93), .A2(Y1_4xDP[6]), .ZN(
        mult_lsb_gf4_mul_0_1_n72) );
  XOR2_X1 mult_lsb_gf4_mul_0_1_U24 ( .A(mult_lsb_gf4_mul_0_1_n74), .B(
        mult_lsb_gf4_mul_0_1_n71), .Z(mult_lsb_gf4_mul_0_1_n73) );
  NOR2_X1 mult_lsb_gf4_mul_0_1_U23 ( .A1(mult_lsb_gf4_mul_0_1_n70), .A2(
        mult_lsb_gf4_mul_0_1_n69), .ZN(mult_lsb_gf4_mul_0_1_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U22 ( .A(n93), .B(n95), .ZN(
        mult_lsb_gf4_mul_0_1_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U21 ( .A(Y1_4xDP[6]), .B(Y1_4xDP[7]), .ZN(
        mult_lsb_gf4_mul_0_1_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U20 ( .A(mult_lsb_gf4_mul_0_1_n68), .B(
        mult_lsb_gf4_mul_0_1_n67), .ZN(mult_lsb_Xi_mul_Yj_1__1_) );
  NAND2_X1 mult_lsb_gf4_mul_0_1_U19 ( .A1(n91), .A2(Y1_4xDP[5]), .ZN(
        mult_lsb_gf4_mul_0_1_n67) );
  XOR2_X1 mult_lsb_gf4_mul_0_1_U18 ( .A(mult_lsb_gf4_mul_0_1_n75), .B(
        mult_lsb_gf4_mul_0_1_n66), .Z(mult_lsb_gf4_mul_0_1_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U17 ( .A(mult_lsb_gf4_mul_0_1_n65), .B(
        mult_lsb_gf4_mul_0_1_n64), .ZN(mult_lsb_gf4_mul_0_1_n75) );
  NAND2_X1 mult_lsb_gf4_mul_0_1_U16 ( .A1(mult_lsb_gf4_mul_0_1_n63), .A2(
        mult_lsb_gf4_mul_0_1_n62), .ZN(mult_lsb_gf4_mul_0_1_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U15 ( .A(mult_lsb_gf4_mul_0_1_n61), .B(
        mult_lsb_gf4_mul_0_1_n60), .ZN(mult_lsb_gf4_mul_0_1_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U14 ( .A(mult_lsb_gf4_mul_0_1_n59), .B(
        mult_lsb_gf4_mul_0_1_n58), .ZN(mult_lsb_gf4_mul_0_1_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U13 ( .A(mult_lsb_gf4_mul_0_1_n57), .B(
        mult_lsb_gf4_mul_0_1_n56), .ZN(mult_lsb_Xi_mul_Yj_1__0_) );
  NAND2_X1 mult_lsb_gf4_mul_0_1_U12 ( .A1(n89), .A2(Y1_4xDP[4]), .ZN(
        mult_lsb_gf4_mul_0_1_n56) );
  XOR2_X1 mult_lsb_gf4_mul_0_1_U11 ( .A(mult_lsb_gf4_mul_0_1_n66), .B(
        mult_lsb_gf4_mul_0_1_n71), .Z(mult_lsb_gf4_mul_0_1_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U10 ( .A(mult_lsb_gf4_mul_0_1_n55), .B(
        mult_lsb_gf4_mul_0_1_n65), .ZN(mult_lsb_gf4_mul_0_1_n71) );
  NOR2_X1 mult_lsb_gf4_mul_0_1_U9 ( .A1(mult_lsb_gf4_mul_0_1_n61), .A2(
        mult_lsb_gf4_mul_0_1_n59), .ZN(mult_lsb_gf4_mul_0_1_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U8 ( .A(n89), .B(n93), .ZN(
        mult_lsb_gf4_mul_0_1_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U7 ( .A(Y1_4xDP[4]), .B(Y1_4xDP[6]), .ZN(
        mult_lsb_gf4_mul_0_1_n61) );
  NAND2_X1 mult_lsb_gf4_mul_0_1_U6 ( .A1(mult_lsb_gf4_mul_0_1_n58), .A2(
        mult_lsb_gf4_mul_0_1_n60), .ZN(mult_lsb_gf4_mul_0_1_n55) );
  XOR2_X1 mult_lsb_gf4_mul_0_1_U5 ( .A(Y1_4xDP[5]), .B(Y1_4xDP[7]), .Z(
        mult_lsb_gf4_mul_0_1_n60) );
  XOR2_X1 mult_lsb_gf4_mul_0_1_U4 ( .A(n91), .B(n95), .Z(
        mult_lsb_gf4_mul_0_1_n58) );
  NOR2_X1 mult_lsb_gf4_mul_0_1_U3 ( .A1(mult_lsb_gf4_mul_0_1_n54), .A2(
        mult_lsb_gf4_mul_0_1_n53), .ZN(mult_lsb_gf4_mul_0_1_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U2 ( .A(n89), .B(n91), .ZN(
        mult_lsb_gf4_mul_0_1_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_0_1_U1 ( .A(Y1_4xDP[4]), .B(Y1_4xDP[5]), .ZN(
        mult_lsb_gf4_mul_0_1_n54) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U29 ( .A(mult_lsb_gf4_mul_0_0_n77), .B(
        mult_lsb_gf4_mul_0_0_n76), .ZN(mult_lsb_FFxDN[3]) );
  NAND2_X1 mult_lsb_gf4_mul_0_0_U28 ( .A1(n95), .A2(Y1_4xDP[3]), .ZN(
        mult_lsb_gf4_mul_0_0_n76) );
  XOR2_X1 mult_lsb_gf4_mul_0_0_U27 ( .A(mult_lsb_gf4_mul_0_0_n75), .B(
        mult_lsb_gf4_mul_0_0_n74), .Z(mult_lsb_gf4_mul_0_0_n77) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U26 ( .A(mult_lsb_gf4_mul_0_0_n73), .B(
        mult_lsb_gf4_mul_0_0_n72), .ZN(mult_lsb_FFxDN[2]) );
  NAND2_X1 mult_lsb_gf4_mul_0_0_U25 ( .A1(n93), .A2(Y1_4xDP[2]), .ZN(
        mult_lsb_gf4_mul_0_0_n72) );
  XOR2_X1 mult_lsb_gf4_mul_0_0_U24 ( .A(mult_lsb_gf4_mul_0_0_n74), .B(
        mult_lsb_gf4_mul_0_0_n71), .Z(mult_lsb_gf4_mul_0_0_n73) );
  NOR2_X1 mult_lsb_gf4_mul_0_0_U23 ( .A1(mult_lsb_gf4_mul_0_0_n70), .A2(
        mult_lsb_gf4_mul_0_0_n69), .ZN(mult_lsb_gf4_mul_0_0_n74) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U22 ( .A(n93), .B(n95), .ZN(
        mult_lsb_gf4_mul_0_0_n69) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U21 ( .A(Y1_4xDP[2]), .B(Y1_4xDP[3]), .ZN(
        mult_lsb_gf4_mul_0_0_n70) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U20 ( .A(mult_lsb_gf4_mul_0_0_n68), .B(
        mult_lsb_gf4_mul_0_0_n67), .ZN(mult_lsb_FFxDN[1]) );
  NAND2_X1 mult_lsb_gf4_mul_0_0_U19 ( .A1(n91), .A2(Y1_4xDP[1]), .ZN(
        mult_lsb_gf4_mul_0_0_n67) );
  XOR2_X1 mult_lsb_gf4_mul_0_0_U18 ( .A(mult_lsb_gf4_mul_0_0_n75), .B(
        mult_lsb_gf4_mul_0_0_n66), .Z(mult_lsb_gf4_mul_0_0_n68) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U17 ( .A(mult_lsb_gf4_mul_0_0_n65), .B(
        mult_lsb_gf4_mul_0_0_n64), .ZN(mult_lsb_gf4_mul_0_0_n75) );
  NAND2_X1 mult_lsb_gf4_mul_0_0_U16 ( .A1(mult_lsb_gf4_mul_0_0_n63), .A2(
        mult_lsb_gf4_mul_0_0_n62), .ZN(mult_lsb_gf4_mul_0_0_n64) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U15 ( .A(mult_lsb_gf4_mul_0_0_n61), .B(
        mult_lsb_gf4_mul_0_0_n60), .ZN(mult_lsb_gf4_mul_0_0_n62) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U14 ( .A(mult_lsb_gf4_mul_0_0_n59), .B(
        mult_lsb_gf4_mul_0_0_n58), .ZN(mult_lsb_gf4_mul_0_0_n63) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U13 ( .A(mult_lsb_gf4_mul_0_0_n57), .B(
        mult_lsb_gf4_mul_0_0_n56), .ZN(mult_lsb_FFxDN[0]) );
  NAND2_X1 mult_lsb_gf4_mul_0_0_U12 ( .A1(n89), .A2(Y1_4xDP[0]), .ZN(
        mult_lsb_gf4_mul_0_0_n56) );
  XOR2_X1 mult_lsb_gf4_mul_0_0_U11 ( .A(mult_lsb_gf4_mul_0_0_n66), .B(
        mult_lsb_gf4_mul_0_0_n71), .Z(mult_lsb_gf4_mul_0_0_n57) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U10 ( .A(mult_lsb_gf4_mul_0_0_n55), .B(
        mult_lsb_gf4_mul_0_0_n65), .ZN(mult_lsb_gf4_mul_0_0_n71) );
  NOR2_X1 mult_lsb_gf4_mul_0_0_U9 ( .A1(mult_lsb_gf4_mul_0_0_n61), .A2(
        mult_lsb_gf4_mul_0_0_n59), .ZN(mult_lsb_gf4_mul_0_0_n65) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U8 ( .A(n89), .B(n93), .ZN(
        mult_lsb_gf4_mul_0_0_n59) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U7 ( .A(Y1_4xDP[0]), .B(Y1_4xDP[2]), .ZN(
        mult_lsb_gf4_mul_0_0_n61) );
  NAND2_X1 mult_lsb_gf4_mul_0_0_U6 ( .A1(mult_lsb_gf4_mul_0_0_n58), .A2(
        mult_lsb_gf4_mul_0_0_n60), .ZN(mult_lsb_gf4_mul_0_0_n55) );
  XOR2_X1 mult_lsb_gf4_mul_0_0_U5 ( .A(Y1_4xDP[1]), .B(Y1_4xDP[3]), .Z(
        mult_lsb_gf4_mul_0_0_n60) );
  XOR2_X1 mult_lsb_gf4_mul_0_0_U4 ( .A(n91), .B(n95), .Z(
        mult_lsb_gf4_mul_0_0_n58) );
  NOR2_X1 mult_lsb_gf4_mul_0_0_U3 ( .A1(mult_lsb_gf4_mul_0_0_n54), .A2(
        mult_lsb_gf4_mul_0_0_n53), .ZN(mult_lsb_gf4_mul_0_0_n66) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U2 ( .A(n89), .B(n91), .ZN(
        mult_lsb_gf4_mul_0_0_n53) );
  XNOR2_X1 mult_lsb_gf4_mul_0_0_U1 ( .A(Y1_4xDP[0]), .B(Y1_4xDP[1]), .ZN(
        mult_lsb_gf4_mul_0_0_n54) );
endmodule

